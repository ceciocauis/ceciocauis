magic
tech sky130A
timestamp 1681049173
<< nwell >>
rect 19000 13700 20500 16200
rect 21100 13700 22600 16200
rect 23200 13700 24700 16200
<< pwell >>
rect 18000 16200 25500 30000
rect 18000 13700 19000 16200
rect 20500 13700 21100 16200
rect 22600 13700 23200 16200
rect 24700 13700 25500 16200
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 19200 27800 20300 27810
rect 19200 26590 20300 26600
rect 21280 27800 22420 27810
rect 21280 26600 21300 27800
rect 22400 26600 22420 27800
rect 21280 26590 22420 26600
rect 23400 27800 24500 27810
rect 23400 26590 24500 26600
rect 18880 16300 24820 16310
rect 18880 13600 18900 16300
rect 24800 13600 24820 16300
rect 18880 13590 24820 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 19100 13810 19120 16100
rect 19280 15000 20220 15010
rect 19280 14000 19300 15000
rect 20200 14000 20220 15000
rect 19280 13990 20220 14000
rect 20380 13810 20400 16100
rect 19100 13800 20400 13810
rect 21200 13810 21220 16100
rect 21380 15000 22320 15010
rect 21380 14000 21400 15000
rect 22300 14000 22320 15000
rect 21380 13990 22320 14000
rect 22480 13810 22500 16100
rect 21200 13800 22500 13810
rect 23300 13810 23320 16100
rect 23480 15000 24420 15010
rect 23480 14000 23500 15000
rect 24400 14000 24420 15000
rect 23480 13990 24420 14000
rect 24580 13810 24600 16100
rect 23300 13800 24600 13810
<< psubdiffcont >>
rect 18220 27810 25280 29790
rect 18220 26590 19200 27810
rect 20300 26590 21280 27810
rect 22420 26590 23400 27810
rect 24500 26590 25280 27810
rect 18220 16310 25280 26590
rect 18220 13590 18880 16310
rect 24820 13590 25280 16310
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 19120 15010 20380 16100
rect 19120 13990 19280 15010
rect 20220 13990 20380 15010
rect 19120 13810 20380 13990
rect 21220 15010 22480 16100
rect 21220 13990 21380 15010
rect 22320 13990 22480 15010
rect 21220 13810 22480 13990
rect 23320 15010 24580 16100
rect 23320 13990 23480 15010
rect 24420 13990 24580 15010
rect 23320 13810 24580 13990
<< pdiode >>
rect 19300 14690 20200 15000
rect 19300 14310 19610 14690
rect 19890 14310 20200 14690
rect 19300 14000 20200 14310
rect 21400 14690 22300 15000
rect 21400 14310 21710 14690
rect 21990 14310 22300 14690
rect 21400 14000 22300 14310
rect 23500 14690 24400 15000
rect 23500 14310 23810 14690
rect 24090 14310 24400 14690
rect 23500 14000 24400 14310
<< ndiode >>
rect 19300 27390 20200 27700
rect 19300 27010 19610 27390
rect 19890 27010 20200 27390
rect 19300 26700 20200 27010
rect 21400 27390 22300 27700
rect 21400 27010 21710 27390
rect 21990 27010 22300 27390
rect 21400 26700 22300 27010
rect 23500 27390 24400 27700
rect 23500 27010 23810 27390
rect 24090 27010 24400 27390
rect 23500 26700 24400 27010
<< pdiodec >>
rect 19610 14310 19890 14690
rect 21710 14310 21990 14690
rect 23810 14310 24090 14690
<< ndiodec >>
rect 19610 27010 19890 27390
rect 21710 27010 21990 27390
rect 23810 27010 24090 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 19190 29790 24510 29990
rect 19200 27500 20300 27810
rect 21280 27790 22420 27810
rect 19200 26900 19500 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20300 27500
rect 19200 26590 20300 26900
rect 21290 27500 22410 27790
rect 21290 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22410 27500
rect 21290 26590 22410 26900
rect 23400 27500 24500 27810
rect 23400 26900 23700 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24500 27500
rect 23400 26590 24500 26900
rect 18890 16300 24810 16310
rect 18890 13600 18900 16300
rect 19000 16190 24700 16200
rect 19000 13710 19010 16190
rect 19190 16100 20310 16190
rect 21290 16100 22410 16190
rect 23390 16100 24510 16190
rect 19280 14800 20220 15010
rect 19280 14200 19500 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20220 14800
rect 19280 13990 20220 14200
rect 21380 14800 22320 15010
rect 21380 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22320 14800
rect 21380 13990 22320 14200
rect 23480 14800 24420 15010
rect 23480 14200 23700 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24420 14800
rect 23480 13990 24420 14200
rect 19190 13710 20310 13810
rect 21290 13710 22410 13810
rect 23390 13710 24510 13810
rect 24690 13710 24700 16190
rect 19000 13700 24700 13710
rect 24800 13600 24810 16300
rect 18890 13590 24810 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 19190 29990
rect 24510 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 16310 19190 29790
rect 19610 27010 19890 27390
rect 20310 26590 21280 27790
rect 21280 26590 21290 27790
rect 21710 27010 21990 27390
rect 22410 26590 22420 27790
rect 22420 26590 23390 27790
rect 23810 27010 24090 27390
rect 20310 16310 21290 26590
rect 22410 16310 23390 26590
rect 24510 16310 25280 29790
rect 18220 13590 18880 16310
rect 18880 13590 18890 16310
rect 19010 16100 19190 16190
rect 20310 16100 21290 16190
rect 22410 16100 23390 16190
rect 24510 16100 24690 16190
rect 19010 13810 19120 16100
rect 19120 13810 19190 16100
rect 19610 14310 19890 14690
rect 20310 13810 20380 16100
rect 20380 13810 21220 16100
rect 21220 13810 21290 16100
rect 21710 14310 21990 14690
rect 22410 13810 22480 16100
rect 22480 13810 23320 16100
rect 23320 13810 23390 16100
rect 23810 14310 24090 14690
rect 24510 13810 24580 16100
rect 24580 13810 24690 16100
rect 19010 13710 19190 13810
rect 20310 13710 21290 13810
rect 22410 13710 23390 13810
rect 24510 13710 24690 13810
rect 24810 13590 24820 16310
rect 24820 13590 25280 16310
rect 18220 11610 19190 13590
rect 24510 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 19200 30000
rect 18000 11610 18010 29990
rect 19190 16310 19200 29990
rect 18890 16300 19200 16310
rect 19300 27900 24400 30000
rect 19300 27690 20200 27900
rect 19300 26710 19310 27690
rect 20190 26710 20200 27690
rect 18890 13600 18900 16300
rect 19000 16190 19200 16200
rect 19000 13710 19010 16190
rect 19190 13710 19200 16190
rect 19000 13700 19200 13710
rect 19300 14990 20200 26710
rect 20300 27790 21300 27800
rect 20300 16310 20310 27790
rect 21290 16310 21300 27790
rect 20300 16300 21300 16310
rect 21400 27690 22300 27900
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 19300 14010 19310 14990
rect 20190 14010 20200 14990
rect 19300 13600 20200 14010
rect 20300 16190 21300 16200
rect 20300 13710 20310 16190
rect 21290 13710 21300 16190
rect 20300 13700 21300 13710
rect 21400 14990 22300 26710
rect 22400 27790 23400 27800
rect 22400 16310 22410 27790
rect 23390 16310 23400 27790
rect 22400 16300 23400 16310
rect 23500 27690 24400 27900
rect 23500 26710 23510 27690
rect 24390 26710 24400 27690
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 21400 13600 22300 14010
rect 22400 16190 23400 16200
rect 22400 13710 22410 16190
rect 23390 13710 23400 16190
rect 22400 13700 23400 13710
rect 23500 14990 24400 26710
rect 24500 29990 25500 30000
rect 24500 16310 24510 29990
rect 24500 16300 24810 16310
rect 23500 14010 23510 14990
rect 24390 14010 24400 14990
rect 23500 13600 24400 14010
rect 24500 16190 24700 16200
rect 24500 13710 24510 16190
rect 24690 13710 24700 16190
rect 24500 13700 24700 13710
rect 24800 13600 24810 16300
rect 18890 13590 19200 13600
rect 19190 11610 19200 13590
rect 18000 11600 19200 11610
rect 19300 11500 24400 13600
rect 24500 13590 24810 13600
rect 24500 11610 24510 13590
rect 25490 11610 25500 29990
rect 24500 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 19190 29990
rect 19310 27390 20190 27690
rect 19310 27010 19610 27390
rect 19610 27010 19890 27390
rect 19890 27010 20190 27390
rect 19310 26710 20190 27010
rect 19010 13710 19190 16190
rect 20310 20910 21290 27790
rect 21410 27390 22290 27690
rect 21410 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22290 27390
rect 21410 26710 22290 27010
rect 19310 14690 20190 14990
rect 19310 14310 19610 14690
rect 19610 14310 19890 14690
rect 19890 14310 20190 14690
rect 19310 14010 20190 14310
rect 20310 13710 21290 16190
rect 22410 20910 23390 27790
rect 23510 27390 24390 27690
rect 23510 27010 23810 27390
rect 23810 27010 24090 27390
rect 24090 27010 24390 27390
rect 23510 26710 24390 27010
rect 21410 14690 22290 14990
rect 21410 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22290 14690
rect 21410 14010 22290 14310
rect 22410 13710 23390 16190
rect 24510 20910 25490 29990
rect 23510 14690 24390 14990
rect 23510 14310 23810 14690
rect 23810 14310 24090 14690
rect 24090 14310 24390 14690
rect 23510 14010 24390 14310
rect 24510 13710 24690 16190
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19190 27800 20310 27810
rect 19190 26600 19200 27800
rect 19300 27690 20200 27700
rect 19300 26710 19310 27690
rect 20190 26710 20200 27690
rect 19300 26700 20200 26710
rect 20300 26600 20310 27800
rect 21290 27800 22410 27810
rect 19190 26590 20310 26600
rect 21290 26600 21300 27800
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 22400 26600 22410 27800
rect 23390 27800 24510 27810
rect 21290 26590 22410 26600
rect 23390 26600 23400 27800
rect 23500 27690 24400 27700
rect 23500 26710 23510 27690
rect 24390 26710 24400 27690
rect 23500 26700 24400 26710
rect 24500 26600 24510 27800
rect 23390 26590 24510 26600
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19190 15100 20310 15110
rect 19190 13900 19200 15100
rect 19300 14990 20200 15000
rect 19300 14010 19310 14990
rect 20190 14010 20200 14990
rect 19300 14000 20200 14010
rect 20300 13900 20310 15100
rect 19190 13890 20310 13900
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 23390 15100 24510 15110
rect 23390 13900 23400 15100
rect 23500 14990 24400 15000
rect 23500 14010 23510 14990
rect 24390 14010 24400 14990
rect 23500 14000 24400 14010
rect 24500 13900 24510 15100
rect 23390 13890 24510 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 19190 29990
rect 19190 27810 24510 29990
rect 19310 26710 20190 27690
rect 20310 27790 21290 27810
rect 19190 20910 20310 26590
rect 20310 20910 21290 27790
rect 21410 26710 22290 27690
rect 22410 27790 23390 27810
rect 21290 20910 22410 26590
rect 22410 20910 23390 27790
rect 23510 26710 24390 27690
rect 23390 20910 24510 26590
rect 24510 20910 25490 29990
rect 18010 16190 25490 20690
rect 18010 13710 19010 16190
rect 19010 13710 19190 16190
rect 19190 15110 20310 16190
rect 19310 14010 20190 14990
rect 19190 13710 20310 13890
rect 20310 13710 21290 16190
rect 21290 15110 22410 16190
rect 21410 14010 22290 14990
rect 21290 13710 22410 13890
rect 22410 13710 23390 16190
rect 23390 15110 24510 16190
rect 23510 14010 24390 14990
rect 23390 13710 24510 13890
rect 24510 13710 24690 16190
rect 24690 13710 25490 16190
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19200 27800 20310 27810
rect 19200 26610 19210 27800
rect 19300 27690 20200 27700
rect 19300 26710 19310 27690
rect 20190 26710 20200 27690
rect 19300 26700 20200 26710
rect 20300 26610 20310 27800
rect 19200 26600 20310 26610
rect 21290 27800 22410 27810
rect 21290 26610 21300 27800
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 22400 26610 22410 27800
rect 21290 26600 22410 26610
rect 23390 27800 24510 27810
rect 23390 26610 23400 27800
rect 23500 27690 24400 27700
rect 23500 26710 23510 27690
rect 24390 26710 24400 27690
rect 23500 26700 24400 26710
rect 24500 26610 24510 27800
rect 23390 26600 24510 26610
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19200 15100 20310 15110
rect 19200 13900 19210 15100
rect 19300 14990 20200 15000
rect 19300 14010 19310 14990
rect 20190 14010 20200 14990
rect 19300 14000 20200 14010
rect 20300 13900 20310 15100
rect 19200 13890 20310 13900
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 23390 15100 24510 15110
rect 23390 13900 23400 15100
rect 23500 14990 24400 15000
rect 23500 14010 23510 14990
rect 24390 14010 24400 14990
rect 23500 14000 24400 14010
rect 24500 13900 24510 15100
rect 23390 13890 24510 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27810 25490 29990
rect 18010 26590 19190 27810
rect 19190 26600 19200 27810
rect 19310 26710 20190 27690
rect 19190 26590 20310 26600
rect 20310 26590 21290 27810
rect 21410 26710 22290 27690
rect 21290 26590 22410 26600
rect 22410 26590 23390 27810
rect 23510 26710 24390 27690
rect 23390 26590 24510 26600
rect 24510 26590 25490 27810
rect 18010 20910 25490 26590
rect 18010 15110 25490 20690
rect 18010 13890 19190 15110
rect 19190 13890 19200 15110
rect 19310 14010 20190 14990
rect 20310 13890 21290 15110
rect 21410 14010 22290 14990
rect 22410 13890 23390 15110
rect 23510 14010 24390 14990
rect 24510 13890 25490 15110
rect 18010 11610 25490 13890
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19200 27800 20310 27810
rect 19200 26610 19210 27800
rect 20300 26610 20310 27800
rect 19200 26600 20310 26610
rect 21290 27800 22410 27810
rect 21290 26610 21300 27800
rect 22400 26610 22410 27800
rect 21290 26600 22410 26610
rect 23390 27800 24510 27810
rect 23390 26610 23400 27800
rect 24500 26610 24510 27800
rect 23390 26600 24510 26610
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19200 15100 20310 15110
rect 19200 13900 19210 15100
rect 20300 13900 20310 15100
rect 19200 13890 20310 13900
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 23390 15100 24510 15110
rect 23390 13900 23400 15100
rect 24500 13900 24510 15100
rect 23390 13890 24510 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 19300 27690 20200 27700
rect 19300 26710 19310 27690
rect 19310 26710 20190 27690
rect 20190 26710 20200 27690
rect 19300 26700 20200 26710
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 21410 26710 22290 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 23500 27690 24400 27700
rect 23500 26710 23510 27690
rect 23510 26710 24390 27690
rect 24390 26710 24400 27690
rect 23500 26700 24400 26710
rect 19300 14990 20200 15000
rect 19300 14010 19310 14990
rect 19310 14010 20190 14990
rect 20190 14010 20200 14990
rect 19300 14000 20200 14010
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 21410 14010 22290 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
rect 23500 14990 24400 15000
rect 23500 14010 23510 14990
rect 23510 14010 24390 14990
rect 24390 14010 24400 14990
rect 23500 14000 24400 14010
<< metal5 >>
rect 19200 27700 24500 27800
rect 19200 26700 19300 27700
rect 20200 26700 21400 27700
rect 22300 26700 23500 27700
rect 24400 26700 24500 27700
rect 19200 15000 24500 26700
rect 19200 14000 19300 15000
rect 20200 14000 21400 15000
rect 22300 14000 23500 15000
rect 24400 14000 24500 15000
rect 19200 13900 24500 14000
<< labels >>
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
<< end >>
