magic
tech sky130A
timestamp 1679025881
<< nwell >>
rect 19000 13700 20500 18700
rect 21100 13700 22600 18700
rect 23200 13700 24700 18700
<< pwell >>
rect 18000 18700 25500 30000
rect 18000 13700 19000 18700
rect 20500 13700 21100 18700
rect 22600 13700 23200 18700
rect 24700 13700 25500 18700
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 18880 18800 24820 18810
rect 18880 13600 18900 18800
rect 24800 13600 24820 18800
rect 18880 13590 24820 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 19100 13810 19120 18600
rect 19500 18100 20000 18200
rect 19500 17700 19600 18100
rect 19900 17700 20000 18100
rect 19500 17600 20000 17700
rect 19500 14700 20000 14800
rect 19500 14300 19600 14700
rect 19900 14300 20000 14700
rect 19500 14200 20000 14300
rect 20380 13810 20400 18600
rect 19100 13800 20400 13810
rect 21200 13810 21220 18600
rect 21600 18100 22100 18200
rect 21600 17700 21700 18100
rect 22000 17700 22100 18100
rect 21600 17600 22100 17700
rect 21600 14700 22100 14800
rect 21600 14300 21700 14700
rect 22000 14300 22100 14700
rect 21600 14200 22100 14300
rect 22480 13810 22500 18600
rect 21200 13800 22500 13810
rect 23300 13810 23320 18600
rect 23700 18100 24200 18200
rect 23700 17700 23800 18100
rect 24100 17700 24200 18100
rect 23700 17600 24200 17700
rect 23700 14700 24200 14800
rect 23700 14300 23800 14700
rect 24100 14300 24200 14700
rect 23700 14200 24200 14300
rect 24580 13810 24600 18600
rect 23300 13800 24600 13810
<< psubdiffcont >>
rect 18220 27500 25280 29790
rect 18220 26900 19500 27500
rect 20000 26900 21600 27500
rect 22100 26900 23700 27500
rect 24200 26900 25280 27500
rect 18220 24100 25280 26900
rect 18220 23500 19500 24100
rect 20000 23500 21600 24100
rect 22100 23500 23700 24100
rect 24200 23500 25280 24100
rect 18220 18810 25280 23500
rect 18220 13590 18880 18810
rect 24820 13590 25280 18810
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 19120 18200 20380 18600
rect 19120 17600 19500 18200
rect 20000 17600 20380 18200
rect 19120 14800 20380 17600
rect 19120 14200 19500 14800
rect 20000 14200 20380 14800
rect 19120 13810 20380 14200
rect 21220 18200 22480 18600
rect 21220 17600 21600 18200
rect 22100 17600 22480 18200
rect 21220 14800 22480 17600
rect 21220 14200 21600 14800
rect 22100 14200 22480 14800
rect 21220 13810 22480 14200
rect 23320 18200 24580 18600
rect 23320 17600 23700 18200
rect 24200 17600 24580 18200
rect 23320 14800 24580 17600
rect 23320 14200 23700 14800
rect 24200 14200 24580 14800
rect 23320 13810 24580 14200
<< pdiode >>
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
<< ndiode >>
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
<< pdiodec >>
rect 19610 17710 19890 18090
rect 19610 14310 19890 14690
rect 21710 17710 21990 18090
rect 21710 14310 21990 14690
rect 23810 17710 24090 18090
rect 23810 14310 24090 14690
<< ndiodec >>
rect 19610 27010 19890 27390
rect 21710 27010 21990 27390
rect 23810 27010 24090 27390
rect 19610 23610 19890 23990
rect 21710 23610 21990 23990
rect 23810 23610 24090 23990
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 19490 29790 24210 29990
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
rect 18890 18800 24810 18810
rect 18890 13600 18900 18800
rect 19000 18690 24700 18700
rect 19000 13710 19010 18690
rect 19490 18600 20010 18690
rect 21590 18600 22110 18690
rect 23690 18600 24210 18690
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 19490 13710 20010 13810
rect 21590 13710 22110 13810
rect 23690 13710 24210 13810
rect 24690 13710 24700 18690
rect 19000 13700 24700 13710
rect 24800 13600 24810 18800
rect 18890 13590 24810 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 19490 29990
rect 24210 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 18810 19490 29790
rect 19610 27010 19890 27390
rect 19610 23610 19890 23990
rect 20010 18810 21590 27790
rect 21710 27010 21990 27390
rect 21710 23610 21990 23990
rect 22110 18810 23690 27790
rect 23810 27010 24090 27390
rect 23810 23610 24090 23990
rect 24210 18810 25280 29790
rect 18220 13590 18880 18810
rect 18880 13590 18890 18810
rect 19010 18600 19490 18690
rect 20010 18600 21590 18690
rect 22110 18600 23690 18690
rect 24210 18600 24690 18690
rect 19010 13810 19120 18600
rect 19120 13810 19490 18600
rect 19610 17710 19890 18090
rect 19610 14310 19890 14690
rect 20010 13810 20380 18600
rect 20380 13810 21220 18600
rect 21220 13810 21590 18600
rect 21710 17710 21990 18090
rect 21710 14310 21990 14690
rect 22110 13810 22480 18600
rect 22480 13810 23320 18600
rect 23320 13810 23690 18600
rect 23810 17710 24090 18090
rect 23810 14310 24090 14690
rect 24210 13810 24580 18600
rect 24580 13810 24690 18600
rect 19010 13710 19490 13810
rect 20010 13710 21590 13810
rect 22110 13710 23690 13810
rect 24210 13710 24690 13810
rect 24810 13590 24820 18810
rect 24820 13590 25280 18810
rect 18220 11610 19490 13590
rect 24210 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 19500 30000
rect 18000 11610 18010 29990
rect 19490 18810 19500 29990
rect 18890 18800 19500 18810
rect 19600 27900 24100 30000
rect 19600 27390 19900 27900
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 23990 19900 27010
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 18890 13600 18900 18800
rect 19000 18690 19500 18700
rect 19000 13710 19010 18690
rect 19490 13710 19500 18690
rect 19000 13700 19500 13710
rect 19600 18090 19900 23610
rect 20000 27790 21600 27800
rect 20000 18810 20010 27790
rect 21590 18810 21600 27790
rect 20000 18800 21600 18810
rect 21700 27390 22000 27900
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 23990 22000 27010
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 14690 19900 17710
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 13600 19900 14310
rect 20000 18690 21600 18700
rect 20000 13710 20010 18690
rect 21590 13710 21600 18690
rect 20000 13700 21600 13710
rect 21700 18090 22000 23610
rect 22100 27790 23700 27800
rect 22100 18810 22110 27790
rect 23690 18810 23700 27790
rect 22100 18800 23700 18810
rect 23800 27390 24100 27900
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 23990 24100 27010
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 14690 22000 17710
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 13600 22000 14310
rect 22100 18690 23700 18700
rect 22100 13710 22110 18690
rect 23690 13710 23700 18690
rect 22100 13700 23700 13710
rect 23800 18090 24100 23610
rect 24200 29990 25500 30000
rect 24200 18810 24210 29990
rect 24200 18800 24810 18810
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 14690 24100 17710
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 13600 24100 14310
rect 24200 18690 24700 18700
rect 24200 13710 24210 18690
rect 24690 13710 24700 18690
rect 24200 13700 24700 13710
rect 24800 13600 24810 18800
rect 18890 13590 19500 13600
rect 19490 11610 19500 13590
rect 18000 11600 19500 11610
rect 19600 11500 24100 13600
rect 24200 13590 24810 13600
rect 24200 11610 24210 13590
rect 25490 11610 25500 29990
rect 24200 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 19490 29990
rect 19610 27010 19890 27390
rect 19610 23610 19890 23990
rect 19010 13710 19490 18690
rect 21710 27010 21990 27390
rect 21710 23610 21990 23990
rect 19610 17710 19890 18090
rect 19610 14310 19890 14690
rect 20010 13710 21590 18690
rect 23810 27010 24090 27390
rect 23810 23610 24090 23990
rect 21710 17710 21990 18090
rect 21710 14310 21990 14690
rect 22110 13710 23690 18690
rect 24210 20910 25490 29990
rect 23810 17710 24090 18090
rect 23810 14310 24090 14690
rect 24210 13710 24690 18690
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19490 27500 20010 27510
rect 19490 26900 19500 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20010 27500
rect 19490 26890 20010 26900
rect 21590 27500 22110 27510
rect 21590 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22110 27500
rect 21590 26890 22110 26900
rect 23690 27500 24210 27510
rect 23690 26900 23700 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24210 27500
rect 23690 26890 24210 26900
rect 19490 24100 20010 24110
rect 19490 23500 19500 24100
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 20000 23500 20010 24100
rect 19490 23490 20010 23500
rect 21590 24100 22110 24110
rect 21590 23500 21600 24100
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 22100 23500 22110 24100
rect 21590 23490 22110 23500
rect 23690 24100 24210 24110
rect 23690 23500 23700 24100
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
rect 24200 23500 24210 24100
rect 23690 23490 24210 23500
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19490 18200 20010 18210
rect 19490 17600 19500 18200
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 20000 17600 20010 18200
rect 19490 17590 20010 17600
rect 19490 14800 20010 14810
rect 19490 14200 19500 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20010 14800
rect 19490 14190 20010 14200
rect 21590 18200 22110 18210
rect 21590 17600 21600 18200
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 22100 17600 22110 18200
rect 21590 17590 22110 17600
rect 21590 14800 22110 14810
rect 21590 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22110 14800
rect 21590 14190 22110 14200
rect 23690 18200 24210 18210
rect 23690 17600 23700 18200
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 24200 17600 24210 18200
rect 23690 17590 24210 17600
rect 23690 14800 24210 14810
rect 23690 14200 23700 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24210 14800
rect 23690 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 19490 29990
rect 19490 27510 24210 29990
rect 19610 27010 19890 27390
rect 20010 26890 21590 27510
rect 21710 27010 21990 27390
rect 22110 26890 23690 27510
rect 23810 27010 24090 27390
rect 19490 24110 24210 26890
rect 19610 23610 19890 23990
rect 20010 23490 21590 24110
rect 21710 23610 21990 23990
rect 22110 23490 23690 24110
rect 23810 23610 24090 23990
rect 19490 20910 24210 23490
rect 24210 20910 25490 29990
rect 18010 18690 25490 20690
rect 18010 13710 19010 18690
rect 19010 13710 19490 18690
rect 19490 18210 20010 18690
rect 19610 17710 19890 18090
rect 19490 14810 20010 17590
rect 19610 14310 19890 14690
rect 19490 13710 20010 14190
rect 20010 13710 21590 18690
rect 21590 18210 22110 18690
rect 21710 17710 21990 18090
rect 21590 14810 22110 17590
rect 21710 14310 21990 14690
rect 21590 13710 22110 14190
rect 22110 13710 23690 18690
rect 23690 18210 24210 18690
rect 23810 17710 24090 18090
rect 23690 14810 24210 17590
rect 23810 14310 24090 14690
rect 23690 13710 24210 14190
rect 24210 13710 24690 18690
rect 24690 13710 25490 18690
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19500 27500 20010 27510
rect 19500 26900 19510 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20010 27500
rect 19500 26890 20010 26900
rect 21600 27500 22110 27510
rect 21600 26900 21610 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22110 27500
rect 21600 26890 22110 26900
rect 23700 27500 24210 27510
rect 23700 26900 23710 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24210 27500
rect 23700 26890 24210 26900
rect 19500 24100 20010 24110
rect 19500 23500 19510 24100
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 20000 23500 20010 24100
rect 19500 23490 20010 23500
rect 21600 24100 22110 24110
rect 21600 23500 21610 24100
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 22100 23500 22110 24100
rect 21600 23490 22110 23500
rect 23700 24100 24210 24110
rect 23700 23500 23710 24100
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
rect 24200 23500 24210 24100
rect 23700 23490 24210 23500
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19500 18200 20010 18210
rect 19500 17600 19510 18200
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 20000 17600 20010 18200
rect 19500 17590 20010 17600
rect 21600 18200 22110 18210
rect 21600 17600 21610 18200
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 22100 17600 22110 18200
rect 21600 17590 22110 17600
rect 23700 18200 24210 18210
rect 23700 17600 23710 18200
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 24200 17600 24210 18200
rect 23700 17590 24210 17600
rect 19500 14800 20010 14810
rect 19500 14200 19510 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20010 14800
rect 19500 14190 20010 14200
rect 21600 14800 22110 14810
rect 21600 14200 21610 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22110 14800
rect 21600 14190 22110 14200
rect 23700 14800 24210 14810
rect 23700 14200 23710 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24210 14800
rect 23700 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27510 25490 29990
rect 18010 26890 19490 27510
rect 19490 26890 19500 27510
rect 19610 27010 19890 27390
rect 20010 26890 21590 27510
rect 21590 26890 21600 27510
rect 21710 27010 21990 27390
rect 22110 26890 23690 27510
rect 23690 26890 23700 27510
rect 23810 27010 24090 27390
rect 24210 26890 25490 27510
rect 18010 24110 25490 26890
rect 18010 23490 19490 24110
rect 19490 23490 19500 24110
rect 19610 23610 19890 23990
rect 20010 23490 21590 24110
rect 21590 23490 21600 24110
rect 21710 23610 21990 23990
rect 22110 23490 23690 24110
rect 23690 23490 23700 24110
rect 23810 23610 24090 23990
rect 24210 23490 25490 24110
rect 18010 20910 25490 23490
rect 18010 18210 25490 20690
rect 18010 17590 19490 18210
rect 19490 17590 19500 18210
rect 19610 17710 19890 18090
rect 20010 17590 21590 18210
rect 21590 17590 21600 18210
rect 21710 17710 21990 18090
rect 22110 17590 23690 18210
rect 23690 17590 23700 18210
rect 23810 17710 24090 18090
rect 24210 17590 25490 18210
rect 18010 14810 25490 17590
rect 18010 14190 19490 14810
rect 19490 14190 19500 14810
rect 19610 14310 19890 14690
rect 20010 14190 21590 14810
rect 21590 14190 21600 14810
rect 21710 14310 21990 14690
rect 22110 14190 23690 14810
rect 23690 14190 23700 14810
rect 23810 14310 24090 14690
rect 24210 14190 25490 14810
rect 18010 11610 25490 14190
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19500 27500 20010 27510
rect 19500 26900 19510 27500
rect 20000 26900 20010 27500
rect 19500 26890 20010 26900
rect 21600 27500 22110 27510
rect 21600 26900 21610 27500
rect 22100 26900 22110 27500
rect 21600 26890 22110 26900
rect 23700 27500 24210 27510
rect 23700 26900 23710 27500
rect 24200 26900 24210 27500
rect 23700 26890 24210 26900
rect 19500 24100 20010 24110
rect 19500 23500 19510 24100
rect 20000 23500 20010 24100
rect 19500 23490 20010 23500
rect 21600 24100 22110 24110
rect 21600 23500 21610 24100
rect 22100 23500 22110 24100
rect 21600 23490 22110 23500
rect 23700 24100 24210 24110
rect 23700 23500 23710 24100
rect 24200 23500 24210 24100
rect 23700 23490 24210 23500
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19500 18200 20010 18210
rect 19500 17600 19510 18200
rect 20000 17600 20010 18200
rect 19500 17590 20010 17600
rect 21600 18200 22110 18210
rect 21600 17600 21610 18200
rect 22100 17600 22110 18200
rect 21600 17590 22110 17600
rect 23700 18200 24210 18210
rect 23700 17600 23710 18200
rect 24200 17600 24210 18200
rect 23700 17590 24210 17600
rect 19500 14800 20010 14810
rect 19500 14200 19510 14800
rect 20000 14200 20010 14800
rect 19500 14190 20010 14200
rect 21600 14800 22110 14810
rect 21600 14200 21610 14800
rect 22100 14200 22110 14800
rect 21600 14190 22110 14200
rect 23700 14800 24210 14810
rect 23700 14200 23710 14800
rect 24200 14200 24210 14800
rect 23700 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19610 27010 19890 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 23810 27010 24090 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19610 23610 19890 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21710 23610 21990 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 23810 23610 24090 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19610 17710 19890 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21710 17710 21990 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 23810 17710 24090 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19610 14310 19890 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 23810 14310 24090 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
<< metal5 >>
rect 19200 27400 24500 27800
rect 19200 27000 19600 27400
rect 19900 27000 21700 27400
rect 22000 27000 23800 27400
rect 24100 27000 24500 27400
rect 19200 24000 24500 27000
rect 19200 23600 19600 24000
rect 19900 23600 21700 24000
rect 22000 23600 23800 24000
rect 24100 23600 24500 24000
rect 19200 18100 24500 23600
rect 19200 17700 19600 18100
rect 19900 17700 21700 18100
rect 22000 17700 23800 18100
rect 24100 17700 24500 18100
rect 19200 14700 24500 17700
rect 19200 14300 19600 14700
rect 19900 14300 21700 14700
rect 22000 14300 23800 14700
rect 24100 14300 24500 14700
rect 19200 13900 24500 14300
<< labels >>
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
<< end >>
