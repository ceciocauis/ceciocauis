* NGSPICE file created from Padtest.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m5_SYR7BF m5_n1000000_200# m5_n1000000_n257# m5_n1000000_n200#
+ SUB
R0 m5_n1000000_n257# m5_n1000000_200# sky130_fd_pr__res_generic_m5 w=10k w=2
C0 m5_n1000000_n257# SUB 406.53fF
C1 m5_n1000000_n200# SUB 126.56fF
C2 m5_n1000000_200# SUB 406.53fF
.ends

.subckt SigPad_6x7_2di vdd vss in
D0 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=2.6e+07 area=4.2e+13
D1 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=2.6e+07 area=4.2e+13
C0 vdd in 378.20fF
C1 in vss 656.38fF
C2 vdd vss 881.61fF
.ends

.subckt Padtest in out vss vdd
XR1 in out R1/m5_n1000000_n200# vss sky130_fd_pr__res_generic_m5_SYR7BF
XSigPad_6x7_2di_0 vdd vss out SigPad_6x7_2di
R0 out.t0 out 0.921
R1 out.t0 out.t1 0.067
R2 out out.t0 0.003
R3 vdd.n0 vdd 0.022
R4 vdd.n1 vdd 0.014
R5 vdd vdd.n6 0.012
R6 vdd.n5 vdd.n0 0.009
R7 vdd.n4 vdd.n3 0.006
R8 vdd.n2 vdd.n1 0.006
R9 vdd.n6 vdd.n5 0.006
R10 vdd.n4 vdd.n2 0.005
R11 vdd.n5 vdd.n4 0.005
R12 vss.n15 vss.n12 10.794
R13 vss.n6 vss.n5 4.461
R14 vss.n19 vss.n18 4.247
R15 vss.n19 vss.n16 2.474
R16 vss.n16 vss.n15 1.066
R17 vss.n18 vss.n17 0.73
R18 vss.n9 vss.n7 0.142
R19 vss.n9 vss.n8 0.134
R20 vss.n2 vss 0.084
R21 vss.n10 vss.n9 0.086
R22 vss.n11 vss.n10 0.052
R23 vss.n23 vss.n22 0.016
R24 vss.n21 vss.n1 0.014
R25 vss vss.n23 0.013
R26 vss.n2 vss 0.012
R27 vss.n3 vss.n2 0.006
R28 vss.n23 vss.n21 0.006
R29 vss.n6 vss.n4 0.006
R30 vss.n20 vss.n19 0.005
R31 vss.n11 vss.n6 0.001
R32 vss.n14 vss.n13 0.001
R33 vss.n15 vss.n14 0.001
R34 vss.n19 vss.n11 0.001
R35 vss.n4 vss.n3 0.001
R36 vss.n1 vss.n0 0.001
R37 vss.n21 vss.n20 0.001
C0 vdd out -1.71fF
C1 out R1/m5_n1000000_n200# 2.13fF
C2 vdd in 13.34fF
C3 vdd R1/m5_n1000000_n200# 12.62fF
C4 out in 1.47fF
C5 vdd.n0 vss 204.39fF $ **FLOATING
C6 vdd.n1 vss 70.64fF $ **FLOATING
C7 vdd.n2 vss 309.07fF $ **FLOATING
C8 vdd.n3 vss 317.82fF $ **FLOATING
C9 vdd.n5 vss 233.62fF $ **FLOATING
C10 vdd.n6 vss 68.59fF $ **FLOATING
C11 out.t1 vss 410.50fF
C12 out.t0 vss 761.88fF
C13 out vss 1305.04fF
C14 vdd vss 961.54fF
C15 R1/m5_n1000000_n200# vss 139.33fF
C16 in vss 842.06fF
.ends

