* NGSPICE file created from Padtest.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m5_SYR7BF m5_n1000000_200# m5_n1000000_n257# m5_n1000000_n200#
+ SUB
R0 m5_n1000000_n257# m5_n1000000_200# sky130_fd_pr__res_generic_m5 w=10k w=2
C0 m5_n1000000_n257# SUB 406.53fF
C1 m5_n1000000_n200# SUB 126.56fF
C2 m5_n1000000_200# SUB 406.53fF
.ends

.subckt SigPad_9x10_6di vdd vss in
D0 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D1 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D2 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D3 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D4 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D5 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
C0 vdd in 791.99fF
C1 in vss 1514.88fF
C2 vdd vss 573.80fF
.ends

.subckt Padtest in out vss vdd
XR1 in out R1/m5_n1000000_n200# vss sky130_fd_pr__res_generic_m5_SYR7BF
XSigPad_9x10_6di_0 vdd vss out SigPad_9x10_6di
R0 out.t1 out 0.36
R1 out.t1 out.n0 0.063
R2 out.n0 out.t2 0.003
R3 out out.t1 0.002
R4 out.n0 out.t0 0.001
R5 vss.n44 vss.n38 142.894
R6 vss.n36 vss.n35 38.939
R7 vss.n28 vss.n27 4.624
R8 vss.n40 vss.n39 2.543
R9 vss.n24 vss.n23 1.323
R10 vss.n24 vss.n18 1.23
R11 vss.n42 vss.n40 0.518
R12 vss.n42 vss.n41 0.419
R13 vss.n11 vss 0.268
R14 vss.n45 vss.n44 0.181
R15 vss.n45 vss.n37 0.178
R16 vss.n44 vss.n43 0.127
R17 vss.n34 vss.n33 0.097
R18 vss.n29 vss.n26 0.086
R19 vss.n22 vss.n21 0.072
R20 vss.n24 vss.n22 0.061
R21 vss.n2 vss.n1 0.059
R22 vss.n3 vss.n0 0.054
R23 vss.n30 vss.n29 0.051
R24 vss.n34 vss.n30 0.05
R25 vss.n29 vss.n28 0.049
R26 vss.n6 vss 0.043
R27 vss.n37 vss.n36 0.033
R28 vss.n43 vss.n42 0.028
R29 vss.n47 vss.n10 0.027
R30 vss.n16 vss.n15 0.027
R31 vss.n8 vss.n6 0.023
R32 vss.n49 vss.n8 0.022
R33 vss.n24 vss.n20 0.02
R34 vss.n5 vss.n4 0.02
R35 vss.n45 vss.n17 0.02
R36 vss.n49 vss.n48 0.009
R37 vss.n12 vss.n11 0.008
R38 vss.n13 vss.n12 0.008
R39 vss.n46 vss.n13 0.008
R40 vss.n48 vss.n47 0.008
R41 vss.n47 vss.n46 0.007
R42 vss.n6 vss.n5 0.006
R43 vss.n45 vss.n25 0.006
R44 vss.n25 vss.n24 0.006
R45 vss.n45 vss.n14 0.006
R46 vss vss.n49 0.004
R47 vss.n46 vss.n45 0.004
R48 vss.n11 vss 0.003
R49 vss.n37 vss.n34 0.003
R50 vss.n3 vss.n2 0.002
R51 vss.n10 vss.n9 0.001
R52 vss.n17 vss.n16 0.001
R53 vss.n32 vss.n31 0.001
R54 vss.n33 vss.n32 0.001
R55 vss.n20 vss.n19 0.001
R56 vss.n5 vss.n3 0.001
R57 vss.n8 vss.n7 0.001
R58 vdd.n25 vdd.n24 5.094
R59 vdd.n2 vdd.n1 2.269
R60 vdd.n18 vdd.n17 1.668
R61 vdd.n34 vdd.n33 1.613
R62 vdd.n34 vdd.n32 0.767
R63 vdd.n35 vdd.n34 0.612
R64 vdd.n17 vdd.n16 0.154
R65 vdd.n4 vdd 0.108
R66 vdd.n31 vdd.n28 0.075
R67 vdd.n11 vdd.n6 0.075
R68 vdd.n3 vdd.n0 0.037
R69 vdd.n23 vdd.n22 0.034
R70 vdd.n31 vdd.n29 0.028
R71 vdd.n31 vdd.n30 0.028
R72 vdd.n39 vdd.n11 0.028
R73 vdd.n11 vdd.n8 0.028
R74 vdd.n11 vdd.n10 0.028
R75 vdd.n40 vdd.n5 0.028
R76 vdd.n5 vdd.n4 0.028
R77 vdd.n38 vdd.n15 0.023
R78 vdd.n8 vdd.n7 0.023
R79 vdd.n38 vdd.n14 0.021
R80 vdd.n10 vdd.n9 0.021
R81 vdd.n13 vdd.n12 0.018
R82 vdd.n40 vdd.n39 0.017
R83 vdd.n3 vdd.n2 0.016
R84 vdd.n35 vdd.n31 0.015
R85 vdd.n25 vdd.n23 0.014
R86 vdd.n39 vdd.n38 0.009
R87 vdd.n20 vdd.n19 0.008
R88 vdd.n38 vdd.n20 0.008
R89 vdd.n37 vdd.n36 0.008
R90 vdd.n4 vdd 0.008
R91 vdd.n27 vdd.n26 0.007
R92 vdd.n37 vdd.n35 0.007
R93 vdd.n20 vdd.n18 0.007
R94 vdd.n38 vdd.n37 0.007
R95 vdd.n38 vdd.n13 0.007
R96 vdd.n12 vdd 0.005
R97 vdd vdd.n40 0.003
R98 vdd.n26 vdd.n25 0.001
R99 vdd.n5 vdd.n3 0.001
R100 vdd.n23 vdd.n21 0.001
R101 vdd.n35 vdd.n27 0.001
C0 R1/m5_n1000000_n200# vdd 12.62fF
C1 in vdd 13.34fF
C2 out R1/m5_n1000000_n200# 2.13fF
C3 out vdd -1.71fF
C4 out in 1.47fF
C5 vdd.n0 vss 47.78fF $ **FLOATING
C6 vdd.n1 vss 3.68fF $ **FLOATING
C7 vdd.n2 vss 45.41fF $ **FLOATING
C8 vdd.n3 vss 9.80fF $ **FLOATING
C9 vdd.n4 vss 26.17fF $ **FLOATING
C10 vdd.n5 vss 13.70fF $ **FLOATING
C11 vdd.n6 vss 16.43fF $ **FLOATING
C12 vdd.n7 vss 29.22fF $ **FLOATING
C13 vdd.n8 vss 24.43fF $ **FLOATING
C14 vdd.n9 vss 16.00fF $ **FLOATING
C15 vdd.n10 vss 16.43fF $ **FLOATING
C16 vdd.n11 vss 9.98fF $ **FLOATING
C17 vdd.n12 vss 49.63fF $ **FLOATING
C18 vdd.n13 vss 55.09fF $ **FLOATING
C19 vdd.n14 vss 34.33fF $ **FLOATING
C20 vdd.n15 vss 36.03fF $ **FLOATING
C21 vdd.n16 vss 3.44fF $ **FLOATING
C22 vdd.n17 vss 9.68fF $ **FLOATING
C23 vdd.n18 vss 78.67fF $ **FLOATING
C24 vdd.n19 vss 103.01fF $ **FLOATING
C25 vdd.n20 vss 36.03fF $ **FLOATING
C26 vdd.n21 vss 34.53fF $ **FLOATING
C27 vdd.n22 vss 49.18fF $ **FLOATING
C28 vdd.n23 vss 12.21fF $ **FLOATING
C29 vdd.n24 vss 4.02fF $ **FLOATING
C30 vdd.n25 vss 59.11fF $ **FLOATING
C31 vdd.n26 vss 12.94fF $ **FLOATING
C32 vdd.n27 vss 34.28fF $ **FLOATING
C33 vdd.n28 vss 15.73fF $ **FLOATING
C34 vdd.n29 vss 32.58fF $ **FLOATING
C35 vdd.n30 vss 15.73fF $ **FLOATING
C36 vdd.n31 vss 9.98fF $ **FLOATING
C37 vdd.n32 vss 12.59fF $ **FLOATING
C38 vdd.n33 vss 32.06fF $ **FLOATING
C39 vdd.n35 vss 33.06fF $ **FLOATING
C40 vdd.n36 vss 104.03fF $ **FLOATING
C41 vdd.n37 vss 34.33fF $ **FLOATING
C42 vdd.n38 vss 110.11fF $ **FLOATING
C43 vdd.n39 vss 56.87fF $ **FLOATING
C44 vdd.n40 vss 44.16fF $ **FLOATING
C45 out.t2 vss 160.48fF
C46 out.t0 vss 844.63fF
C47 out.n0 vss 46.52fF $ **FLOATING
C48 out.t1 vss 1706.01fF
C49 out vss 1850.54fF
C50 vdd vss 591.43fF
C51 R1/m5_n1000000_n200# vss 139.33fF
C52 in vss 842.06fF
.ends

