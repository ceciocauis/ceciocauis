* NGSPICE file created from Padtest.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m5_SYR7BF m5_n1000000_200# m5_n1000000_n257# m5_n1000000_n200#
+ SUB
R0 m5_n1000000_n257# m5_n1000000_200# sky130_fd_pr__res_generic_m5 w=10k w=2
C0 m5_n1000000_n257# SUB 406.53fF
C1 m5_n1000000_n200# SUB 126.56fF
C2 m5_n1000000_200# SUB 406.53fF
.ends

.subckt SigPad_3x4_4di vdd vss in
D0 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=1.4e+07 area=1.2e+13
D1 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=1.4e+07 area=1.2e+13
D2 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=1.4e+07 area=1.2e+13
D3 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=1.4e+07 area=1.2e+13
C0 in vdd 506.40fF
C1 in vss 989.31fF
C2 vdd vss 730.71fF
.ends

.subckt Padtest in out vss vdd
XR1 in out R1/m5_n1000000_n200# vss sky130_fd_pr__res_generic_m5_SYR7BF
XSigPad_3x4_4di_0 vdd vss out SigPad_3x4_4di
R0 out.t2 out 0.537
R1 out.t0 out.n0 0.386
R2 out.t2 out.n1 0.069
R3 out out.t2 0.003
R4 out.n1 out.t1 0.003
R5 out.n1 out.t0 0.001
R6 vss vss.n11 14.004
R7 vss vss.n10 7.072
R8 vss.n10 vss.n9 5.951
R9 vss.n4 vss.n3 0.255
R10 vss.n0 vss 0.216
R11 vss.n6 vss.n4 0.21
R12 vss.n1 vss 0.178
R13 vss vss.n15 0.128
R14 vss.n15 vss.n12 0.086
R15 vss.n8 vss.n7 0.058
R16 vss.n7 vss.n6 0.033
R17 vss vss.n2 0.011
R18 vss.n2 vss.n0 0.01
R19 vss vss.n8 0.006
R20 vss.n2 vss.n1 0.005
R21 vss.n0 vss 0.004
R22 vss.n6 vss.n5 0.001
R23 vss.n15 vss.n14 0.001
R24 vss.n14 vss.n13 0.001
R25 vdd vdd.n10 0.094
R26 vdd.n10 vdd.n9 0.034
R27 vdd.n9 vdd 0.034
R28 vdd.n2 vdd 0.015
R29 vdd.n4 vdd.n3 0.012
R30 vdd.n8 vdd.n0 0.01
R31 vdd.n10 vdd.n8 0.01
R32 vdd.n8 vdd.n4 0.007
R33 vdd.n8 vdd.n5 0.005
R34 vdd.n0 vdd 0.004
R35 vdd.n3 vdd.n1 0.001
R36 vdd.n3 vdd.n2 0.001
R37 vdd.n8 vdd.n7 0.001
R38 vdd.n7 vdd.n6 0.001
C0 out R1/m5_n1000000_n200# 2.13fF
C1 out in 1.47fF
C2 R1/m5_n1000000_n200# vdd 12.62fF
C3 in vdd 13.34fF
C4 out vdd -1.71fF
C5 vdd.n0 vss 59.14fF $ **FLOATING
C6 vdd.n1 vss 18.79fF $ **FLOATING
C7 vdd.n2 vss 176.26fF $ **FLOATING
C8 vdd.n3 vss 450.23fF $ **FLOATING
C9 vdd.n4 vss 98.18fF $ **FLOATING
C10 vdd.n5 vss 45.81fF $ **FLOATING
C11 vdd.n6 vss 39.28fF $ **FLOATING
C12 vdd.n7 vss 47.28fF $ **FLOATING
C13 vdd.n8 vss 43.10fF $ **FLOATING
C14 vdd.n9 vss 29.96fF $ **FLOATING
C15 vdd.n10 vss 16.92fF $ **FLOATING
C16 out.t1 vss -17.11fF
C17 out.t0 vss 94.21fF
C18 out.n1 vss 554.75fF $ **FLOATING
C19 out.t2 vss 1121.97fF
C20 out vss 1517.65fF
C21 vdd vss 967.13fF
C22 R1/m5_n1000000_n200# vss 139.33fF
C23 in vss 842.06fF
.ends

