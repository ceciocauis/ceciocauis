magic
tech sky130A
timestamp 1679065267
<< nwell >>
rect 21100 13700 22600 15300
<< pwell >>
rect 18000 15300 25500 30000
rect 18000 13700 21100 15300
rect 22600 13700 25500 15300
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 20980 15400 22720 15410
rect 20980 13600 21000 15400
rect 22700 13600 22720 15400
rect 20980 13590 22720 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 21200 13810 21220 15200
rect 21600 14700 22100 14800
rect 21600 14300 21700 14700
rect 22000 14300 22100 14700
rect 21600 14200 22100 14300
rect 22480 13810 22500 15200
rect 21200 13800 22500 13810
<< psubdiffcont >>
rect 18220 27500 25280 29790
rect 18220 26900 21600 27500
rect 22100 26900 25280 27500
rect 18220 15410 25280 26900
rect 18220 13590 20980 15410
rect 22720 13590 25280 15410
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 21220 14800 22480 15200
rect 21220 14200 21600 14800
rect 22100 14200 22480 14800
rect 21220 13810 22480 14200
<< pdiode >>
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
<< ndiode >>
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
<< pdiodec >>
rect 21710 14310 21990 14690
<< ndiodec >>
rect 21710 27010 21990 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 21590 29790 22110 29990
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 20990 15400 22710 15410
rect 20990 13600 21000 15400
rect 21100 15290 22600 15300
rect 21100 13710 21110 15290
rect 21590 15200 22110 15290
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 21590 13710 22110 13810
rect 22590 13710 22600 15290
rect 21100 13700 22600 13710
rect 22700 13600 22710 15400
rect 20990 13590 22710 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 21590 29990
rect 22110 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 15410 21590 29790
rect 21710 27010 21990 27390
rect 22110 15410 25280 29790
rect 18220 13590 20980 15410
rect 20980 13590 20990 15410
rect 21110 15200 21590 15290
rect 22110 15200 22590 15290
rect 21110 13810 21220 15200
rect 21220 13810 21590 15200
rect 21710 14310 21990 14690
rect 22110 13810 22480 15200
rect 22480 13810 22590 15200
rect 21110 13710 21590 13810
rect 22110 13710 22590 13810
rect 22710 13590 22720 15410
rect 22720 13590 25280 15410
rect 18220 11610 21590 13590
rect 22110 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 21600 30000
rect 18000 11610 18010 29990
rect 21590 15410 21600 29990
rect 20990 15400 21600 15410
rect 21700 27390 22000 30000
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 20990 13600 21000 15400
rect 21100 15290 21600 15300
rect 21100 13710 21110 15290
rect 21590 13710 21600 15290
rect 21100 13700 21600 13710
rect 21700 14690 22000 27010
rect 22100 29990 25500 30000
rect 22100 15410 22110 29990
rect 22100 15400 22710 15410
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 20990 13590 21600 13600
rect 21590 11610 21600 13590
rect 18000 11600 21600 11610
rect 21700 11500 22000 14310
rect 22100 15290 22600 15300
rect 22100 13710 22110 15290
rect 22590 13710 22600 15290
rect 22100 13700 22600 13710
rect 22700 13600 22710 15400
rect 22100 13590 22710 13600
rect 22100 11610 22110 13590
rect 25490 11610 25500 29990
rect 22100 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 21590 29990
rect 21710 27010 21990 27390
rect 21110 13710 21590 15290
rect 22110 20910 25490 29990
rect 21710 14310 21990 14690
rect 22110 13710 22590 15290
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21590 27500 22110 27510
rect 21590 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22110 27500
rect 21590 26890 22110 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21590 14800 22110 14810
rect 21590 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22110 14800
rect 21590 14190 22110 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 21590 29990
rect 21590 27510 22110 29990
rect 21710 27010 21990 27390
rect 21590 20910 22110 26890
rect 22110 20910 25490 29990
rect 18010 15290 25490 20690
rect 18010 13710 21110 15290
rect 21110 13710 21590 15290
rect 21590 14810 22110 15290
rect 21710 14310 21990 14690
rect 21590 13710 22110 14190
rect 22110 13710 22590 15290
rect 22590 13710 25490 15290
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21600 27500 22110 27510
rect 21600 26900 21610 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22110 27500
rect 21600 26890 22110 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21600 14800 22110 14810
rect 21600 14200 21610 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22110 14800
rect 21600 14190 22110 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27510 25490 29990
rect 18010 26890 21590 27510
rect 21590 26890 21600 27510
rect 21710 27010 21990 27390
rect 22110 26890 25490 27510
rect 18010 20910 25490 26890
rect 18010 14810 25490 20690
rect 18010 14190 21590 14810
rect 21590 14190 21600 14810
rect 21710 14310 21990 14690
rect 22110 14190 25490 14810
rect 18010 11610 25490 14190
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21600 27500 22110 27510
rect 21600 26900 21610 27500
rect 22100 26900 22110 27500
rect 21600 26890 22110 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21600 14800 22110 14810
rect 21600 14200 21610 14800
rect 22100 14200 22110 14800
rect 21600 14190 22110 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
<< metal5 >>
rect 19200 27400 24500 27800
rect 19200 27000 21700 27400
rect 22000 27000 24500 27400
rect 19200 14700 24500 27000
rect 19200 14300 21700 14700
rect 22000 14300 24500 14700
rect 19200 13900 24500 14300
<< labels >>
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
<< end >>
