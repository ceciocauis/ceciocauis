* NGSPICE file created from Padtest.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m5_SYR7BF m5_n1000000_200# m5_n1000000_n257# m5_n1000000_n200#
+ SUB
R0 m5_n1000000_n257# m5_n1000000_200# sky130_fd_pr__res_generic_m5 w=10k w=2
C0 m5_n1000000_n257# SUB 406.53fF
C1 m5_n1000000_n200# SUB 126.56fF
C2 m5_n1000000_200# SUB 406.53fF
.ends

.subckt SigPad_9x10_12di vdd vss in
D0 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D1 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D2 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D3 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D4 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D5 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D6 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
D7 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D8 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D9 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D10 vss in sky130_fd_pr__diode_pw2nd_05v5 pj=3.8e+07 area=9e+13
D11 in vdd sky130_fd_pr__diode_pd2nw_05v5 pj=3.8e+07 area=9e+13
C0 in vdd 860.22fF
C1 in vss 1408.79fF
C2 vdd vss 593.08fF
.ends

.subckt Padtest in out vss vdd
XR1 in out R1/m5_n1000000_n200# vss sky130_fd_pr__res_generic_m5_SYR7BF
XSigPad_9x10_12di_0 vdd vss out SigPad_9x10_12di
R0 out.t2 out 0.36
R1 out.t3 out.n0 0.047
R2 out.t3 out.n3 0.032
R3 out.t2 out.n4 0.018
R4 out.n2 out.t0 0.018
R5 out.n1 out.t5 0.003
R6 out.n3 out.t1 0.002
R7 out.n3 out.t6 0.002
R8 out out.t2 0.002
R9 out.n4 out.t4 0.001
R10 out.t6 out.n2 0.001
R11 out.t0 out.n1 0.001
R12 out.n4 out.t3 0.001
R13 vss.n0 vss.n66 147.75
R14 vss.n64 vss.n56 24.625
R15 vss.n51 vss.n50 12.232
R16 vss.n64 vss.n30 10.559
R17 vss.n54 vss.n53 10.444
R18 vss.n68 vss.n67 9.956
R19 vss.n61 vss.n60 2.319
R20 vss.n0 vss.n65 1.772
R21 vss.n70 vss.n69 1.725
R22 vss.n63 vss.n62 1.699
R23 vss.n55 vss.n54 1.23
R24 vss.n53 vss.n52 0.985
R25 vss.n59 vss.n58 0.59
R26 vss.n64 vss.n59 0.545
R27 vss.n69 vss.n68 0.466
R28 vss.n59 vss.n57 0.409
R29 vss.n75 vss 0.268
R30 vss.n64 vss.n63 0.205
R31 vss.n65 vss.n64 0.142
R32 vss.n53 vss.n51 0.117
R33 vss.n19 vss 0.108
R34 vss.n64 vss.n55 0.096
R35 vss.n47 vss.n33 0.067
R36 vss.n6 vss.n5 0.059
R37 vss.n32 vss.n31 0.059
R38 vss.n65 vss.n29 0.059
R39 vss.n40 vss.n39 0.057
R40 vss.n45 vss.n44 0.057
R41 vss.n7 vss.n3 0.054
R42 vss.n11 vss 0.043
R43 vss.n20 vss.n14 0.036
R44 vss.n62 vss.n61 0.036
R45 vss.n46 vss.n45 0.034
R46 vss.n75 vss.n20 0.028
R47 vss.n20 vss.n19 0.028
R48 vss.n43 vss.n37 0.028
R49 vss.n73 vss.n24 0.028
R50 vss.n12 vss.n11 0.027
R51 vss.n75 vss.n12 0.027
R52 vss.n73 vss.n22 0.027
R53 vss.n11 vss.n10 0.027
R54 vss.n48 vss.n32 0.024
R55 vss.n35 vss.n34 0.024
R56 vss.n11 vss.n2 0.023
R57 vss.n48 vss.n47 0.023
R58 vss.n47 vss.n35 0.023
R59 vss.n42 vss.n38 0.023
R60 vss.n17 vss.n16 0.022
R61 vss.n27 vss.n26 0.022
R62 vss.n6 vss.n4 0.022
R63 vss.n75 vss.n74 0.022
R64 vss.n74 vss.n73 0.022
R65 vss.n73 vss.n72 0.022
R66 vss.n14 vss.n13 0.022
R67 vss.n45 vss.n43 0.021
R68 vss.n20 vss.n18 0.021
R69 vss.n71 vss.n0 0.02
R70 vss.n9 vss.n8 0.02
R71 vss.n71 vss.n25 0.02
R72 vss.n43 vss.n42 0.019
R73 vss.n24 vss.n23 0.019
R74 vss.n35 vss 0.012
R75 vss.n0 vss.n70 0.01
R76 vss vss.n75 0.008
R77 vss.n19 vss 0.008
R78 vss.n11 vss.n9 0.006
R79 vss.n2 vss.n1 0.004
R80 vss.n72 vss.n71 0.002
R81 vss.n41 vss.n40 0.002
R82 vss.n28 vss.n27 0.002
R83 vss.n7 vss.n6 0.002
R84 vss.n22 vss.n21 0.001
R85 vss.n18 vss.n17 0.001
R86 vss.n37 vss.n36 0.001
R87 vss.n49 vss.n48 0.001
R88 vss.n71 vss.n28 0.001
R89 vss.n18 vss.n15 0.001
R90 vss.n55 vss.n49 0.001
R91 vss.n9 vss.n7 0.001
R92 vss.n47 vss.n46 0.001
R93 vss.n42 vss.n41 0.001
R94 vdd.n24 vdd 0.268
R95 vdd.n13 vdd 0.108
R96 vdd.n9 vdd.n8 0.059
R97 vdd.n11 vdd 0.043
R98 vdd.n12 vdd.n6 0.036
R99 vdd.n15 vdd.n14 0.036
R100 vdd.n24 vdd.n16 0.028
R101 vdd.n16 vdd.n13 0.028
R102 vdd.n12 vdd.n11 0.027
R103 vdd.n24 vdd.n12 0.027
R104 vdd.n22 vdd.n17 0.027
R105 vdd.n12 vdd.n5 0.027
R106 vdd.n22 vdd.n21 0.024
R107 vdd.n9 vdd.n7 0.022
R108 vdd.n24 vdd.n23 0.022
R109 vdd.n23 vdd.n22 0.022
R110 vdd.n3 vdd.n0 11.099
R111 vdd.n0 vdd 0.012
R112 vdd.n3 vdd.n2 0.01
R113 vdd vdd.n24 0.008
R114 vdd.n13 vdd 0.008
R115 vdd.n11 vdd.n10 0.006
R116 vdd.n4 vdd.n3 0.005
R117 vdd.n4 vdd.n1 0.004
R118 vdd.n21 vdd.n18 0.002
R119 vdd.n10 vdd.n9 0.002
R120 vdd.n5 vdd.n4 0.002
R121 vdd.n21 vdd.n20 0.001
R122 vdd.n16 vdd.n15 0.001
R123 vdd.n20 vdd.n19 0.001
C0 out R1/m5_n1000000_n200# 2.13fF
C1 out vdd -1.71fF
C2 vdd in 13.34fF
C3 out in 1.47fF
C4 vdd R1/m5_n1000000_n200# 12.62fF
C5 vdd.n0 vss 503.71fF $ **FLOATING
C6 vdd.n1 vss 8.58fF $ **FLOATING
C7 vdd.n2 vss 21.67fF $ **FLOATING
C8 vdd.n3 vss 505.56fF $ **FLOATING
C9 vdd.n5 vss 16.23fF $ **FLOATING
C10 vdd.n6 vss 42.44fF $ **FLOATING
C11 vdd.n7 vss 15.55fF $ **FLOATING
C12 vdd.n8 vss 15.27fF $ **FLOATING
C13 vdd.n9 vss 14.62fF $ **FLOATING
C14 vdd.n10 vss 84.88fF $ **FLOATING
C15 vdd.n11 vss 180.64fF $ **FLOATING
C16 vdd.n12 vss 23.50fF $ **FLOATING
C17 vdd.n13 vss 25.00fF $ **FLOATING
C18 vdd.n14 vss 45.42fF $ **FLOATING
C19 vdd.n15 vss 10.03fF $ **FLOATING
C20 vdd.n16 vss 13.52fF $ **FLOATING
C21 vdd.n17 vss 10.38fF $ **FLOATING
C22 vdd.n18 vss 15.26fF $ **FLOATING
C23 vdd.n19 vss 6.07fF $ **FLOATING
C24 vdd.n20 vss 13.41fF $ **FLOATING
C25 vdd.n21 vss 6.60fF $ **FLOATING
C26 vdd.n22 vss 17.60fF $ **FLOATING
C27 vdd.n23 vss 13.41fF $ **FLOATING
C28 vdd.n24 vss 29.20fF $ **FLOATING
C29 out.t4 vss 34.29fF
C30 out.n0 vss 40.79fF $ **FLOATING
C31 out.t1 vss 329.91fF
C32 out.t5 vss 105.76fF
C33 out.n1 vss 15.64fF $ **FLOATING
C34 out.t0 vss 260.20fF
C35 out.n2 vss 67.34fF $ **FLOATING
C36 out.t6 vss 178.92fF
C37 out.n3 vss 89.85fF $ **FLOATING
C38 out.t3 vss 612.45fF
C39 out.n4 vss 7.94fF $ **FLOATING
C40 out.t2 vss 969.17fF
C41 out vss 1751.95fF
C42 vdd vss 432.05fF
C43 R1/m5_n1000000_n200# vss 139.33fF
C44 in vss 842.06fF
.ends

