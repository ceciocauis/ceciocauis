magic
tech sky130A
timestamp 1681048457
<< nwell >>
rect 19000 13700 20500 16200
rect 21100 13700 22600 16200
rect 23200 13700 24700 16200
<< pwell >>
rect 18000 16200 25500 30000
rect 18000 13700 19000 16200
rect 20500 13700 21100 16200
rect 22600 13700 23200 16200
rect 24700 13700 25500 16200
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 19350 27650 20150 27660
rect 19350 26740 20150 26750
rect 21450 27650 22250 27660
rect 21450 26740 22250 26750
rect 23550 27650 24350 27660
rect 23550 26740 24350 26750
rect 18880 16300 24820 16310
rect 18880 13600 18900 16300
rect 24800 13600 24820 16300
rect 18880 13590 24820 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 19100 13810 19120 16100
rect 19430 14850 20070 14860
rect 19430 14150 19450 14850
rect 20050 14150 20070 14850
rect 19430 14140 20070 14150
rect 20380 13810 20400 16100
rect 19100 13800 20400 13810
rect 21200 13810 21220 16100
rect 21530 14850 22170 14860
rect 21530 14150 21550 14850
rect 22150 14150 22170 14850
rect 21530 14140 22170 14150
rect 22480 13810 22500 16100
rect 21200 13800 22500 13810
rect 23300 13810 23320 16100
rect 23630 14850 24270 14860
rect 23630 14150 23650 14850
rect 24250 14150 24270 14850
rect 23630 14140 24270 14150
rect 24580 13810 24600 16100
rect 23300 13800 24600 13810
<< psubdiffcont >>
rect 18220 27660 25280 29790
rect 18220 26740 19350 27660
rect 20150 26740 21450 27660
rect 22250 26740 23550 27660
rect 24350 26740 25280 27660
rect 18220 16310 25280 26740
rect 18220 13590 18880 16310
rect 24820 13590 25280 16310
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 19120 14860 20380 16100
rect 19120 14140 19430 14860
rect 20070 14140 20380 14860
rect 19120 13810 20380 14140
rect 21220 14860 22480 16100
rect 21220 14140 21530 14860
rect 22170 14140 22480 14860
rect 21220 13810 22480 14140
rect 23320 14860 24580 16100
rect 23320 14140 23630 14860
rect 24270 14140 24580 14860
rect 23320 13810 24580 14140
<< pdiode >>
rect 19450 14690 20050 14850
rect 19450 14310 19610 14690
rect 19890 14310 20050 14690
rect 19450 14150 20050 14310
rect 21550 14690 22150 14850
rect 21550 14310 21710 14690
rect 21990 14310 22150 14690
rect 21550 14150 22150 14310
rect 23650 14690 24250 14850
rect 23650 14310 23810 14690
rect 24090 14310 24250 14690
rect 23650 14150 24250 14310
<< ndiode >>
rect 19450 27390 20050 27550
rect 19450 27010 19610 27390
rect 19890 27010 20050 27390
rect 19450 26850 20050 27010
rect 21550 27390 22150 27550
rect 21550 27010 21710 27390
rect 21990 27010 22150 27390
rect 21550 26850 22150 27010
rect 23650 27390 24250 27550
rect 23650 27010 23810 27390
rect 24090 27010 24250 27390
rect 23650 26850 24250 27010
<< pdiodec >>
rect 19610 14310 19890 14690
rect 21710 14310 21990 14690
rect 23810 14310 24090 14690
<< ndiodec >>
rect 19610 27010 19890 27390
rect 21710 27010 21990 27390
rect 23810 27010 24090 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 19340 29790 24360 29990
rect 19350 27500 20150 27660
rect 19350 26900 19500 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20150 27500
rect 19350 26740 20150 26900
rect 21450 27500 22250 27660
rect 21450 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22250 27500
rect 21450 26740 22250 26900
rect 23550 27500 24350 27660
rect 23550 26900 23700 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24350 27500
rect 23550 26740 24350 26900
rect 18890 16300 24810 16310
rect 18890 13600 18900 16300
rect 19000 16190 24700 16200
rect 19000 13710 19010 16190
rect 19340 16100 20160 16190
rect 21440 16100 22260 16190
rect 23540 16100 24360 16190
rect 19430 14800 20070 14860
rect 19430 14200 19500 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20070 14800
rect 19430 14140 20070 14200
rect 21530 14800 22170 14860
rect 21530 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22170 14800
rect 21530 14140 22170 14200
rect 23630 14800 24270 14860
rect 23630 14200 23700 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24270 14800
rect 23630 14140 24270 14200
rect 19340 13710 20160 13810
rect 21440 13710 22260 13810
rect 23540 13710 24360 13810
rect 24690 13710 24700 16190
rect 19000 13700 24700 13710
rect 24800 13600 24810 16300
rect 18890 13590 24810 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 19340 29990
rect 24360 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 16310 19340 29790
rect 19610 27010 19890 27390
rect 20160 16310 21440 27790
rect 21710 27010 21990 27390
rect 22260 16310 23540 27790
rect 23810 27010 24090 27390
rect 24360 16310 25280 29790
rect 18220 13590 18880 16310
rect 18880 13590 18890 16310
rect 19010 16100 19340 16190
rect 20160 16100 21440 16190
rect 22260 16100 23540 16190
rect 24360 16100 24690 16190
rect 19010 13810 19120 16100
rect 19120 13810 19340 16100
rect 19610 14310 19890 14690
rect 20160 13810 20380 16100
rect 20380 13810 21220 16100
rect 21220 13810 21440 16100
rect 21710 14310 21990 14690
rect 22260 13810 22480 16100
rect 22480 13810 23320 16100
rect 23320 13810 23540 16100
rect 23810 14310 24090 14690
rect 24360 13810 24580 16100
rect 24580 13810 24690 16100
rect 19010 13710 19340 13810
rect 20160 13710 21440 13810
rect 22260 13710 23540 13810
rect 24360 13710 24690 13810
rect 24810 13590 24820 16310
rect 24820 13590 25280 16310
rect 18220 11610 19340 13590
rect 24360 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 19350 30000
rect 18000 11610 18010 29990
rect 19340 16310 19350 29990
rect 18890 16300 19350 16310
rect 19450 27900 24250 30000
rect 19450 27540 20050 27900
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 18890 13600 18900 16300
rect 19000 16190 19350 16200
rect 19000 13710 19010 16190
rect 19340 13710 19350 16190
rect 19000 13700 19350 13710
rect 19450 14840 20050 26860
rect 20150 27790 21450 27800
rect 20150 16310 20160 27790
rect 21440 16310 21450 27790
rect 20150 16300 21450 16310
rect 21550 27540 22150 27900
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 13600 20050 14160
rect 20150 16190 21450 16200
rect 20150 13710 20160 16190
rect 21440 13710 21450 16190
rect 20150 13700 21450 13710
rect 21550 14840 22150 26860
rect 22250 27790 23550 27800
rect 22250 16310 22260 27790
rect 23540 16310 23550 27790
rect 22250 16300 23550 16310
rect 23650 27540 24250 27900
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 13600 22150 14160
rect 22250 16190 23550 16200
rect 22250 13710 22260 16190
rect 23540 13710 23550 16190
rect 22250 13700 23550 13710
rect 23650 14840 24250 26860
rect 24350 29990 25500 30000
rect 24350 16310 24360 29990
rect 24350 16300 24810 16310
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 13600 24250 14160
rect 24350 16190 24700 16200
rect 24350 13710 24360 16190
rect 24690 13710 24700 16190
rect 24350 13700 24700 13710
rect 24800 13600 24810 16300
rect 18890 13590 19350 13600
rect 19340 11610 19350 13590
rect 18000 11600 19350 11610
rect 19450 11500 24250 13600
rect 24350 13590 24810 13600
rect 24350 11610 24360 13590
rect 25490 11610 25500 29990
rect 24350 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 19340 29990
rect 19460 27390 20040 27540
rect 19460 27010 19610 27390
rect 19610 27010 19890 27390
rect 19890 27010 20040 27390
rect 19460 26860 20040 27010
rect 19010 13710 19340 16190
rect 20160 20910 21440 27790
rect 21560 27390 22140 27540
rect 21560 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22140 27390
rect 21560 26860 22140 27010
rect 19460 14690 20040 14840
rect 19460 14310 19610 14690
rect 19610 14310 19890 14690
rect 19890 14310 20040 14690
rect 19460 14160 20040 14310
rect 20160 13710 21440 16190
rect 22260 20910 23540 27790
rect 23660 27390 24240 27540
rect 23660 27010 23810 27390
rect 23810 27010 24090 27390
rect 24090 27010 24240 27390
rect 23660 26860 24240 27010
rect 21560 14690 22140 14840
rect 21560 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22140 14690
rect 21560 14160 22140 14310
rect 22260 13710 23540 16190
rect 24360 20910 25490 29990
rect 23660 14690 24240 14840
rect 23660 14310 23810 14690
rect 23810 14310 24090 14690
rect 24090 14310 24240 14690
rect 23660 14160 24240 14310
rect 24360 13710 24690 16190
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19340 27650 20160 27660
rect 19340 26750 19350 27650
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 20150 26750 20160 27650
rect 19340 26740 20160 26750
rect 21440 27650 22260 27660
rect 21440 26750 21450 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21440 26740 22260 26750
rect 23540 27650 24360 27660
rect 23540 26750 23550 27650
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 24350 26750 24360 27650
rect 23540 26740 24360 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19340 14950 20160 14960
rect 19340 14050 19350 14950
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 20150 14050 20160 14950
rect 19340 14040 20160 14050
rect 21440 14950 22260 14960
rect 21440 14050 21450 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21440 14040 22260 14050
rect 23540 14950 24360 14960
rect 23540 14050 23550 14950
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
rect 24350 14050 24360 14950
rect 23540 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 19340 29990
rect 19340 27790 24360 29990
rect 19340 27660 20160 27790
rect 19460 26860 20040 27540
rect 19340 20910 20160 26740
rect 20160 20910 21440 27790
rect 21440 27660 22260 27790
rect 21560 26860 22140 27540
rect 21440 20910 22260 26740
rect 22260 20910 23540 27790
rect 23540 27660 24360 27790
rect 23660 26860 24240 27540
rect 23540 20910 24360 26740
rect 24360 20910 25490 29990
rect 18010 16190 25490 20690
rect 18010 13710 19010 16190
rect 19010 13710 19340 16190
rect 19340 14960 20160 16190
rect 19460 14160 20040 14840
rect 19340 13710 20160 14040
rect 20160 13710 21440 16190
rect 21440 14960 22260 16190
rect 21560 14160 22140 14840
rect 21440 13710 22260 14040
rect 22260 13710 23540 16190
rect 23540 14960 24360 16190
rect 23660 14160 24240 14840
rect 23540 13710 24360 14040
rect 24360 13710 24690 16190
rect 24690 13710 25490 16190
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19350 27650 20160 27660
rect 19350 26750 19360 27650
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 20150 26750 20160 27650
rect 19350 26740 20160 26750
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 23550 27650 24360 27660
rect 23550 26750 23560 27650
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 24350 26750 24360 27650
rect 23550 26740 24360 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19350 14950 20160 14960
rect 19350 14050 19360 14950
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 20150 14050 20160 14950
rect 19350 14040 20160 14050
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 23550 14950 24360 14960
rect 23550 14050 23560 14950
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
rect 24350 14050 24360 14950
rect 23550 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27660 25490 29990
rect 18010 26740 19340 27660
rect 19340 26740 19350 27660
rect 19460 26860 20040 27540
rect 20160 26740 21440 27660
rect 21440 26740 21450 27660
rect 21560 26860 22140 27540
rect 22260 26740 23540 27660
rect 23540 26740 23550 27660
rect 23660 26860 24240 27540
rect 24360 26740 25490 27660
rect 18010 20910 25490 26740
rect 18010 14960 25490 20690
rect 18010 14040 19340 14960
rect 19340 14040 19350 14960
rect 19460 14160 20040 14840
rect 20160 14040 21440 14960
rect 21440 14040 21450 14960
rect 21560 14160 22140 14840
rect 22260 14040 23540 14960
rect 23540 14040 23550 14960
rect 23660 14160 24240 14840
rect 24360 14040 25490 14960
rect 18010 11610 25490 14040
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19350 27650 20160 27660
rect 19350 26750 19360 27650
rect 20150 26750 20160 27650
rect 19350 26740 20160 26750
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 23550 27650 24360 27660
rect 23550 26750 23560 27650
rect 24350 26750 24360 27650
rect 23550 26740 24360 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19350 14950 20160 14960
rect 19350 14050 19360 14950
rect 20150 14050 20160 14950
rect 19350 14040 20160 14050
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 23550 14950 24360 14960
rect 23550 14050 23560 14950
rect 24350 14050 24360 14950
rect 23550 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 19460 26860 20040 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 21560 26860 22140 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 23660 26860 24240 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 19460 14160 20040 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 21560 14160 22140 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 23660 14160 24240 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
<< metal5 >>
rect 19200 27550 24500 27800
rect 19200 26850 19450 27550
rect 20050 26850 21550 27550
rect 22150 26850 23650 27550
rect 24250 26850 24500 27550
rect 19200 14850 24500 26850
rect 19200 14150 19450 14850
rect 20050 14150 21550 14850
rect 22150 14150 23650 14850
rect 24250 14150 24500 14850
rect 19200 13900 24500 14150
<< labels >>
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
<< end >>
