magic
tech sky130A
timestamp 1679092491
<< nwell >>
rect 19000 13700 20500 18700
rect 21100 13700 22600 18700
rect 23200 13700 24700 18700
<< pwell >>
rect 18000 18700 25500 30000
rect 18000 13700 19000 18700
rect 20500 13700 21100 18700
rect 22600 13700 23200 18700
rect 24700 13700 25500 18700
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 19350 27650 20150 27660
rect 19350 26740 20150 26750
rect 21450 27650 22250 27660
rect 21450 26740 22250 26750
rect 23550 27650 24350 27660
rect 23550 26740 24350 26750
rect 19350 24250 20150 24260
rect 19350 23340 20150 23350
rect 21450 24250 22250 24260
rect 21450 23340 22250 23350
rect 23550 24250 24350 24260
rect 23550 23340 24350 23350
rect 18880 18800 24820 18810
rect 18880 13600 18900 18800
rect 24800 13600 24820 18800
rect 18880 13590 24820 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 19100 13810 19120 18600
rect 19430 18250 20070 18260
rect 19430 17550 19450 18250
rect 20050 17550 20070 18250
rect 19430 17540 20070 17550
rect 19430 14850 20070 14860
rect 19430 14150 19450 14850
rect 20050 14150 20070 14850
rect 19430 14140 20070 14150
rect 20380 13810 20400 18600
rect 19100 13800 20400 13810
rect 21200 13810 21220 18600
rect 21530 18250 22170 18260
rect 21530 17550 21550 18250
rect 22150 17550 22170 18250
rect 21530 17540 22170 17550
rect 21530 14850 22170 14860
rect 21530 14150 21550 14850
rect 22150 14150 22170 14850
rect 21530 14140 22170 14150
rect 22480 13810 22500 18600
rect 21200 13800 22500 13810
rect 23300 13810 23320 18600
rect 23630 18250 24270 18260
rect 23630 17550 23650 18250
rect 24250 17550 24270 18250
rect 23630 17540 24270 17550
rect 23630 14850 24270 14860
rect 23630 14150 23650 14850
rect 24250 14150 24270 14850
rect 23630 14140 24270 14150
rect 24580 13810 24600 18600
rect 23300 13800 24600 13810
<< psubdiffcont >>
rect 18220 27660 25280 29790
rect 18220 26740 19350 27660
rect 20150 26740 21450 27660
rect 22250 26740 23550 27660
rect 24350 26740 25280 27660
rect 18220 24260 25280 26740
rect 18220 23340 19350 24260
rect 20150 23340 21450 24260
rect 22250 23340 23550 24260
rect 24350 23340 25280 24260
rect 18220 18810 25280 23340
rect 18220 13590 18880 18810
rect 24820 13590 25280 18810
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 19120 18260 20380 18600
rect 19120 17540 19430 18260
rect 20070 17540 20380 18260
rect 19120 14860 20380 17540
rect 19120 14140 19430 14860
rect 20070 14140 20380 14860
rect 19120 13810 20380 14140
rect 21220 18260 22480 18600
rect 21220 17540 21530 18260
rect 22170 17540 22480 18260
rect 21220 14860 22480 17540
rect 21220 14140 21530 14860
rect 22170 14140 22480 14860
rect 21220 13810 22480 14140
rect 23320 18260 24580 18600
rect 23320 17540 23630 18260
rect 24270 17540 24580 18260
rect 23320 14860 24580 17540
rect 23320 14140 23630 14860
rect 24270 14140 24580 14860
rect 23320 13810 24580 14140
<< pdiode >>
rect 19450 18090 20050 18250
rect 19450 17710 19610 18090
rect 19890 17710 20050 18090
rect 19450 17550 20050 17710
rect 19450 14690 20050 14850
rect 19450 14310 19610 14690
rect 19890 14310 20050 14690
rect 19450 14150 20050 14310
rect 21550 18090 22150 18250
rect 21550 17710 21710 18090
rect 21990 17710 22150 18090
rect 21550 17550 22150 17710
rect 21550 14690 22150 14850
rect 21550 14310 21710 14690
rect 21990 14310 22150 14690
rect 21550 14150 22150 14310
rect 23650 18090 24250 18250
rect 23650 17710 23810 18090
rect 24090 17710 24250 18090
rect 23650 17550 24250 17710
rect 23650 14690 24250 14850
rect 23650 14310 23810 14690
rect 24090 14310 24250 14690
rect 23650 14150 24250 14310
<< ndiode >>
rect 19450 27390 20050 27550
rect 19450 27010 19610 27390
rect 19890 27010 20050 27390
rect 19450 26850 20050 27010
rect 21550 27390 22150 27550
rect 21550 27010 21710 27390
rect 21990 27010 22150 27390
rect 21550 26850 22150 27010
rect 23650 27390 24250 27550
rect 23650 27010 23810 27390
rect 24090 27010 24250 27390
rect 23650 26850 24250 27010
rect 19450 23990 20050 24150
rect 19450 23610 19610 23990
rect 19890 23610 20050 23990
rect 19450 23450 20050 23610
rect 21550 23990 22150 24150
rect 21550 23610 21710 23990
rect 21990 23610 22150 23990
rect 21550 23450 22150 23610
rect 23650 23990 24250 24150
rect 23650 23610 23810 23990
rect 24090 23610 24250 23990
rect 23650 23450 24250 23610
<< pdiodec >>
rect 19610 17710 19890 18090
rect 19610 14310 19890 14690
rect 21710 17710 21990 18090
rect 21710 14310 21990 14690
rect 23810 17710 24090 18090
rect 23810 14310 24090 14690
<< ndiodec >>
rect 19610 27010 19890 27390
rect 21710 27010 21990 27390
rect 23810 27010 24090 27390
rect 19610 23610 19890 23990
rect 21710 23610 21990 23990
rect 23810 23610 24090 23990
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 19340 29790 24360 29990
rect 19350 27500 20150 27660
rect 19350 26900 19500 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20150 27500
rect 19350 26740 20150 26900
rect 19350 24100 20150 24260
rect 19350 23500 19500 24100
rect 19600 23990 19900 24000
rect 19600 23610 19610 23990
rect 19890 23610 19900 23990
rect 19600 23600 19900 23610
rect 20000 23500 20150 24100
rect 19350 23340 20150 23500
rect 21450 27500 22250 27660
rect 21450 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22250 27500
rect 21450 26740 22250 26900
rect 21450 24100 22250 24260
rect 21450 23500 21600 24100
rect 21700 23990 22000 24000
rect 21700 23610 21710 23990
rect 21990 23610 22000 23990
rect 21700 23600 22000 23610
rect 22100 23500 22250 24100
rect 21450 23340 22250 23500
rect 23550 27500 24350 27660
rect 23550 26900 23700 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24350 27500
rect 23550 26740 24350 26900
rect 23550 24100 24350 24260
rect 23550 23500 23700 24100
rect 23800 23990 24100 24000
rect 23800 23610 23810 23990
rect 24090 23610 24100 23990
rect 23800 23600 24100 23610
rect 24200 23500 24350 24100
rect 23550 23340 24350 23500
rect 18890 18800 24810 18810
rect 18890 13600 18900 18800
rect 19000 18690 24700 18700
rect 19000 13710 19010 18690
rect 19340 18600 20160 18690
rect 21440 18600 22260 18690
rect 23540 18600 24360 18690
rect 19430 18200 20070 18260
rect 19430 17600 19500 18200
rect 19600 18090 19900 18100
rect 19600 17710 19610 18090
rect 19890 17710 19900 18090
rect 19600 17700 19900 17710
rect 20000 17600 20070 18200
rect 19430 17540 20070 17600
rect 19430 14800 20070 14860
rect 19430 14200 19500 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20070 14800
rect 19430 14140 20070 14200
rect 21530 18200 22170 18260
rect 21530 17600 21600 18200
rect 21700 18090 22000 18100
rect 21700 17710 21710 18090
rect 21990 17710 22000 18090
rect 21700 17700 22000 17710
rect 22100 17600 22170 18200
rect 21530 17540 22170 17600
rect 21530 14800 22170 14860
rect 21530 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22170 14800
rect 21530 14140 22170 14200
rect 23630 18200 24270 18260
rect 23630 17600 23700 18200
rect 23800 18090 24100 18100
rect 23800 17710 23810 18090
rect 24090 17710 24100 18090
rect 23800 17700 24100 17710
rect 24200 17600 24270 18200
rect 23630 17540 24270 17600
rect 23630 14800 24270 14860
rect 23630 14200 23700 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24270 14800
rect 23630 14140 24270 14200
rect 19340 13710 20160 13810
rect 21440 13710 22260 13810
rect 23540 13710 24360 13810
rect 24690 13710 24700 18690
rect 19000 13700 24700 13710
rect 24800 13600 24810 18800
rect 18890 13590 24810 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 19340 29990
rect 24360 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 18810 19340 29790
rect 19610 27010 19890 27390
rect 19610 23610 19890 23990
rect 20160 18810 21440 27790
rect 21710 27010 21990 27390
rect 21710 23610 21990 23990
rect 22260 18810 23540 27790
rect 23810 27010 24090 27390
rect 23810 23610 24090 23990
rect 24360 18810 25280 29790
rect 18220 13590 18880 18810
rect 18880 13590 18890 18810
rect 19010 18600 19340 18690
rect 20160 18600 21440 18690
rect 22260 18600 23540 18690
rect 24360 18600 24690 18690
rect 19010 13810 19120 18600
rect 19120 13810 19340 18600
rect 19610 17710 19890 18090
rect 19610 14310 19890 14690
rect 20160 13810 20380 18600
rect 20380 13810 21220 18600
rect 21220 13810 21440 18600
rect 21710 17710 21990 18090
rect 21710 14310 21990 14690
rect 22260 13810 22480 18600
rect 22480 13810 23320 18600
rect 23320 13810 23540 18600
rect 23810 17710 24090 18090
rect 23810 14310 24090 14690
rect 24360 13810 24580 18600
rect 24580 13810 24690 18600
rect 19010 13710 19340 13810
rect 20160 13710 21440 13810
rect 22260 13710 23540 13810
rect 24360 13710 24690 13810
rect 24810 13590 24820 18810
rect 24820 13590 25280 18810
rect 18220 11610 19340 13590
rect 24360 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 19350 30000
rect 18000 11610 18010 29990
rect 19340 18810 19350 29990
rect 18890 18800 19350 18810
rect 19450 27900 24250 30000
rect 19450 27540 20050 27900
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 19450 24140 20050 26860
rect 19450 23460 19460 24140
rect 20040 23460 20050 24140
rect 18890 13600 18900 18800
rect 19000 18690 19350 18700
rect 19000 13710 19010 18690
rect 19340 13710 19350 18690
rect 19000 13700 19350 13710
rect 19450 18240 20050 23460
rect 20150 27790 21450 27800
rect 20150 18810 20160 27790
rect 21440 18810 21450 27790
rect 20150 18800 21450 18810
rect 21550 27540 22150 27900
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 24140 22150 26860
rect 21550 23460 21560 24140
rect 22140 23460 22150 24140
rect 19450 17560 19460 18240
rect 20040 17560 20050 18240
rect 19450 14840 20050 17560
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 13600 20050 14160
rect 20150 18690 21450 18700
rect 20150 13710 20160 18690
rect 21440 13710 21450 18690
rect 20150 13700 21450 13710
rect 21550 18240 22150 23460
rect 22250 27790 23550 27800
rect 22250 18810 22260 27790
rect 23540 18810 23550 27790
rect 22250 18800 23550 18810
rect 23650 27540 24250 27900
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 23650 24140 24250 26860
rect 23650 23460 23660 24140
rect 24240 23460 24250 24140
rect 21550 17560 21560 18240
rect 22140 17560 22150 18240
rect 21550 14840 22150 17560
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 13600 22150 14160
rect 22250 18690 23550 18700
rect 22250 13710 22260 18690
rect 23540 13710 23550 18690
rect 22250 13700 23550 13710
rect 23650 18240 24250 23460
rect 24350 29990 25500 30000
rect 24350 18810 24360 29990
rect 24350 18800 24810 18810
rect 23650 17560 23660 18240
rect 24240 17560 24250 18240
rect 23650 14840 24250 17560
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 13600 24250 14160
rect 24350 18690 24700 18700
rect 24350 13710 24360 18690
rect 24690 13710 24700 18690
rect 24350 13700 24700 13710
rect 24800 13600 24810 18800
rect 18890 13590 19350 13600
rect 19340 11610 19350 13590
rect 18000 11600 19350 11610
rect 19450 11500 24250 13600
rect 24350 13590 24810 13600
rect 24350 11610 24360 13590
rect 25490 11610 25500 29990
rect 24350 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 19340 29990
rect 19460 27390 20040 27540
rect 19460 27010 19610 27390
rect 19610 27010 19890 27390
rect 19890 27010 20040 27390
rect 19460 26860 20040 27010
rect 19460 23990 20040 24140
rect 19460 23610 19610 23990
rect 19610 23610 19890 23990
rect 19890 23610 20040 23990
rect 19460 23460 20040 23610
rect 19010 13710 19340 18690
rect 20160 20910 21440 27790
rect 21560 27390 22140 27540
rect 21560 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22140 27390
rect 21560 26860 22140 27010
rect 21560 23990 22140 24140
rect 21560 23610 21710 23990
rect 21710 23610 21990 23990
rect 21990 23610 22140 23990
rect 21560 23460 22140 23610
rect 19460 18090 20040 18240
rect 19460 17710 19610 18090
rect 19610 17710 19890 18090
rect 19890 17710 20040 18090
rect 19460 17560 20040 17710
rect 19460 14690 20040 14840
rect 19460 14310 19610 14690
rect 19610 14310 19890 14690
rect 19890 14310 20040 14690
rect 19460 14160 20040 14310
rect 20160 13710 21440 18690
rect 22260 20910 23540 27790
rect 23660 27390 24240 27540
rect 23660 27010 23810 27390
rect 23810 27010 24090 27390
rect 24090 27010 24240 27390
rect 23660 26860 24240 27010
rect 23660 23990 24240 24140
rect 23660 23610 23810 23990
rect 23810 23610 24090 23990
rect 24090 23610 24240 23990
rect 23660 23460 24240 23610
rect 21560 18090 22140 18240
rect 21560 17710 21710 18090
rect 21710 17710 21990 18090
rect 21990 17710 22140 18090
rect 21560 17560 22140 17710
rect 21560 14690 22140 14840
rect 21560 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22140 14690
rect 21560 14160 22140 14310
rect 22260 13710 23540 18690
rect 24360 20910 25490 29990
rect 23660 18090 24240 18240
rect 23660 17710 23810 18090
rect 23810 17710 24090 18090
rect 24090 17710 24240 18090
rect 23660 17560 24240 17710
rect 23660 14690 24240 14840
rect 23660 14310 23810 14690
rect 23810 14310 24090 14690
rect 24090 14310 24240 14690
rect 23660 14160 24240 14310
rect 24360 13710 24690 18690
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19340 27650 20160 27660
rect 19340 26750 19350 27650
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 20150 26750 20160 27650
rect 19340 26740 20160 26750
rect 19340 24250 20160 24260
rect 19340 23350 19350 24250
rect 19450 24140 20050 24150
rect 19450 23460 19460 24140
rect 20040 23460 20050 24140
rect 19450 23450 20050 23460
rect 20150 23350 20160 24250
rect 19340 23340 20160 23350
rect 21440 27650 22260 27660
rect 21440 26750 21450 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21440 26740 22260 26750
rect 21440 24250 22260 24260
rect 21440 23350 21450 24250
rect 21550 24140 22150 24150
rect 21550 23460 21560 24140
rect 22140 23460 22150 24140
rect 21550 23450 22150 23460
rect 22250 23350 22260 24250
rect 21440 23340 22260 23350
rect 23540 27650 24360 27660
rect 23540 26750 23550 27650
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 24350 26750 24360 27650
rect 23540 26740 24360 26750
rect 23540 24250 24360 24260
rect 23540 23350 23550 24250
rect 23650 24140 24250 24150
rect 23650 23460 23660 24140
rect 24240 23460 24250 24140
rect 23650 23450 24250 23460
rect 24350 23350 24360 24250
rect 23540 23340 24360 23350
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19340 18350 20160 18360
rect 19340 17450 19350 18350
rect 19450 18240 20050 18250
rect 19450 17560 19460 18240
rect 20040 17560 20050 18240
rect 19450 17550 20050 17560
rect 20150 17450 20160 18350
rect 19340 17440 20160 17450
rect 19340 14950 20160 14960
rect 19340 14050 19350 14950
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 20150 14050 20160 14950
rect 19340 14040 20160 14050
rect 21440 18350 22260 18360
rect 21440 17450 21450 18350
rect 21550 18240 22150 18250
rect 21550 17560 21560 18240
rect 22140 17560 22150 18240
rect 21550 17550 22150 17560
rect 22250 17450 22260 18350
rect 21440 17440 22260 17450
rect 21440 14950 22260 14960
rect 21440 14050 21450 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21440 14040 22260 14050
rect 23540 18350 24360 18360
rect 23540 17450 23550 18350
rect 23650 18240 24250 18250
rect 23650 17560 23660 18240
rect 24240 17560 24250 18240
rect 23650 17550 24250 17560
rect 24350 17450 24360 18350
rect 23540 17440 24360 17450
rect 23540 14950 24360 14960
rect 23540 14050 23550 14950
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
rect 24350 14050 24360 14950
rect 23540 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 19340 29990
rect 19340 27790 24360 29990
rect 19340 27660 20160 27790
rect 19460 26860 20040 27540
rect 19340 24260 20160 26740
rect 19460 23460 20040 24140
rect 19340 20910 20160 23340
rect 20160 20910 21440 27790
rect 21440 27660 22260 27790
rect 21560 26860 22140 27540
rect 21440 24260 22260 26740
rect 21560 23460 22140 24140
rect 21440 20910 22260 23340
rect 22260 20910 23540 27790
rect 23540 27660 24360 27790
rect 23660 26860 24240 27540
rect 23540 24260 24360 26740
rect 23660 23460 24240 24140
rect 23540 20910 24360 23340
rect 24360 20910 25490 29990
rect 18010 18690 25490 20690
rect 18010 13710 19010 18690
rect 19010 13710 19340 18690
rect 19340 18360 20160 18690
rect 19460 17560 20040 18240
rect 19340 14960 20160 17440
rect 19460 14160 20040 14840
rect 19340 13710 20160 14040
rect 20160 13710 21440 18690
rect 21440 18360 22260 18690
rect 21560 17560 22140 18240
rect 21440 14960 22260 17440
rect 21560 14160 22140 14840
rect 21440 13710 22260 14040
rect 22260 13710 23540 18690
rect 23540 18360 24360 18690
rect 23660 17560 24240 18240
rect 23540 14960 24360 17440
rect 23660 14160 24240 14840
rect 23540 13710 24360 14040
rect 24360 13710 24690 18690
rect 24690 13710 25490 18690
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19350 27650 20160 27660
rect 19350 26750 19360 27650
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 20150 26750 20160 27650
rect 19350 26740 20160 26750
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 23550 27650 24360 27660
rect 23550 26750 23560 27650
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 24350 26750 24360 27650
rect 23550 26740 24360 26750
rect 19350 24250 20160 24260
rect 19350 23350 19360 24250
rect 19450 24140 20050 24150
rect 19450 23460 19460 24140
rect 20040 23460 20050 24140
rect 19450 23450 20050 23460
rect 20150 23350 20160 24250
rect 19350 23340 20160 23350
rect 21450 24250 22260 24260
rect 21450 23350 21460 24250
rect 21550 24140 22150 24150
rect 21550 23460 21560 24140
rect 22140 23460 22150 24140
rect 21550 23450 22150 23460
rect 22250 23350 22260 24250
rect 21450 23340 22260 23350
rect 23550 24250 24360 24260
rect 23550 23350 23560 24250
rect 23650 24140 24250 24150
rect 23650 23460 23660 24140
rect 24240 23460 24250 24140
rect 23650 23450 24250 23460
rect 24350 23350 24360 24250
rect 23550 23340 24360 23350
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19350 18350 20160 18360
rect 19350 17450 19360 18350
rect 19450 18240 20050 18250
rect 19450 17560 19460 18240
rect 20040 17560 20050 18240
rect 19450 17550 20050 17560
rect 20150 17450 20160 18350
rect 19350 17440 20160 17450
rect 21450 18350 22260 18360
rect 21450 17450 21460 18350
rect 21550 18240 22150 18250
rect 21550 17560 21560 18240
rect 22140 17560 22150 18240
rect 21550 17550 22150 17560
rect 22250 17450 22260 18350
rect 21450 17440 22260 17450
rect 23550 18350 24360 18360
rect 23550 17450 23560 18350
rect 23650 18240 24250 18250
rect 23650 17560 23660 18240
rect 24240 17560 24250 18240
rect 23650 17550 24250 17560
rect 24350 17450 24360 18350
rect 23550 17440 24360 17450
rect 19350 14950 20160 14960
rect 19350 14050 19360 14950
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 20150 14050 20160 14950
rect 19350 14040 20160 14050
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 23550 14950 24360 14960
rect 23550 14050 23560 14950
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
rect 24350 14050 24360 14950
rect 23550 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27660 25490 29990
rect 18010 26740 19340 27660
rect 19340 26740 19350 27660
rect 19460 26860 20040 27540
rect 20160 26740 21440 27660
rect 21440 26740 21450 27660
rect 21560 26860 22140 27540
rect 22260 26740 23540 27660
rect 23540 26740 23550 27660
rect 23660 26860 24240 27540
rect 24360 26740 25490 27660
rect 18010 24260 25490 26740
rect 18010 23340 19340 24260
rect 19340 23340 19350 24260
rect 19460 23460 20040 24140
rect 20160 23340 21440 24260
rect 21440 23340 21450 24260
rect 21560 23460 22140 24140
rect 22260 23340 23540 24260
rect 23540 23340 23550 24260
rect 23660 23460 24240 24140
rect 24360 23340 25490 24260
rect 18010 20910 25490 23340
rect 18010 18360 25490 20690
rect 18010 17440 19340 18360
rect 19340 17440 19350 18360
rect 19460 17560 20040 18240
rect 20160 17440 21440 18360
rect 21440 17440 21450 18360
rect 21560 17560 22140 18240
rect 22260 17440 23540 18360
rect 23540 17440 23550 18360
rect 23660 17560 24240 18240
rect 24360 17440 25490 18360
rect 18010 14960 25490 17440
rect 18010 14040 19340 14960
rect 19340 14040 19350 14960
rect 19460 14160 20040 14840
rect 20160 14040 21440 14960
rect 21440 14040 21450 14960
rect 21560 14160 22140 14840
rect 22260 14040 23540 14960
rect 23540 14040 23550 14960
rect 23660 14160 24240 14840
rect 24360 14040 25490 14960
rect 18010 11610 25490 14040
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19350 27650 20160 27660
rect 19350 26750 19360 27650
rect 20150 26750 20160 27650
rect 19350 26740 20160 26750
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 23550 27650 24360 27660
rect 23550 26750 23560 27650
rect 24350 26750 24360 27650
rect 23550 26740 24360 26750
rect 19350 24250 20160 24260
rect 19350 23350 19360 24250
rect 20150 23350 20160 24250
rect 19350 23340 20160 23350
rect 21450 24250 22260 24260
rect 21450 23350 21460 24250
rect 22250 23350 22260 24250
rect 21450 23340 22260 23350
rect 23550 24250 24360 24260
rect 23550 23350 23560 24250
rect 24350 23350 24360 24250
rect 23550 23340 24360 23350
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19350 18350 20160 18360
rect 19350 17450 19360 18350
rect 20150 17450 20160 18350
rect 19350 17440 20160 17450
rect 21450 18350 22260 18360
rect 21450 17450 21460 18350
rect 22250 17450 22260 18350
rect 21450 17440 22260 17450
rect 23550 18350 24360 18360
rect 23550 17450 23560 18350
rect 24350 17450 24360 18350
rect 23550 17440 24360 17450
rect 19350 14950 20160 14960
rect 19350 14050 19360 14950
rect 20150 14050 20160 14950
rect 19350 14040 20160 14050
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 23550 14950 24360 14960
rect 23550 14050 23560 14950
rect 24350 14050 24360 14950
rect 23550 14040 24360 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 19450 27540 20050 27550
rect 19450 26860 19460 27540
rect 19460 26860 20040 27540
rect 20040 26860 20050 27540
rect 19450 26850 20050 26860
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 21560 26860 22140 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 23650 27540 24250 27550
rect 23650 26860 23660 27540
rect 23660 26860 24240 27540
rect 24240 26860 24250 27540
rect 23650 26850 24250 26860
rect 19450 24140 20050 24150
rect 19450 23460 19460 24140
rect 19460 23460 20040 24140
rect 20040 23460 20050 24140
rect 19450 23450 20050 23460
rect 21550 24140 22150 24150
rect 21550 23460 21560 24140
rect 21560 23460 22140 24140
rect 22140 23460 22150 24140
rect 21550 23450 22150 23460
rect 23650 24140 24250 24150
rect 23650 23460 23660 24140
rect 23660 23460 24240 24140
rect 24240 23460 24250 24140
rect 23650 23450 24250 23460
rect 19450 18240 20050 18250
rect 19450 17560 19460 18240
rect 19460 17560 20040 18240
rect 20040 17560 20050 18240
rect 19450 17550 20050 17560
rect 21550 18240 22150 18250
rect 21550 17560 21560 18240
rect 21560 17560 22140 18240
rect 22140 17560 22150 18240
rect 21550 17550 22150 17560
rect 23650 18240 24250 18250
rect 23650 17560 23660 18240
rect 23660 17560 24240 18240
rect 24240 17560 24250 18240
rect 23650 17550 24250 17560
rect 19450 14840 20050 14850
rect 19450 14160 19460 14840
rect 19460 14160 20040 14840
rect 20040 14160 20050 14840
rect 19450 14150 20050 14160
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 21560 14160 22140 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 23650 14840 24250 14850
rect 23650 14160 23660 14840
rect 23660 14160 24240 14840
rect 24240 14160 24250 14840
rect 23650 14150 24250 14160
<< metal5 >>
rect 19200 27550 24500 27800
rect 19200 26850 19450 27550
rect 20050 26850 21550 27550
rect 22150 26850 23650 27550
rect 24250 26850 24500 27550
rect 19200 24150 24500 26850
rect 19200 23450 19450 24150
rect 20050 23450 21550 24150
rect 22150 23450 23650 24150
rect 24250 23450 24500 24150
rect 19200 18250 24500 23450
rect 19200 17550 19450 18250
rect 20050 17550 21550 18250
rect 22150 17550 23650 18250
rect 24250 17550 24500 18250
rect 19200 14850 24500 17550
rect 19200 14150 19450 14850
rect 20050 14150 21550 14850
rect 22150 14150 23650 14850
rect 24250 14150 24500 14850
rect 19200 13900 24500 14150
<< labels >>
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
<< end >>
