magic
tech sky130A
timestamp 1679069139
<< nwell >>
rect 19000 13700 20500 15300
rect 23200 13700 24700 15300
<< pwell >>
rect 18000 15300 25500 30000
rect 18000 13700 19000 15300
rect 20500 13700 23200 15300
rect 24700 13700 25500 15300
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 18880 15400 24820 15410
rect 18880 13600 18900 15400
rect 24800 13600 24820 15400
rect 18880 13590 24820 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 19100 13810 19120 15200
rect 19500 14700 20000 14800
rect 19500 14300 19600 14700
rect 19900 14300 20000 14700
rect 19500 14200 20000 14300
rect 20380 13810 20400 15200
rect 19100 13800 20400 13810
rect 23300 13810 23320 15200
rect 23700 14700 24200 14800
rect 23700 14300 23800 14700
rect 24100 14300 24200 14700
rect 23700 14200 24200 14300
rect 24580 13810 24600 15200
rect 23300 13800 24600 13810
<< psubdiffcont >>
rect 18220 27500 25280 29790
rect 18220 26900 19500 27500
rect 20000 26900 23700 27500
rect 24200 26900 25280 27500
rect 18220 15410 25280 26900
rect 18220 13590 18880 15410
rect 24820 13590 25280 15410
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 19120 14800 20380 15200
rect 19120 14200 19500 14800
rect 20000 14200 20380 14800
rect 19120 13810 20380 14200
rect 23320 14800 24580 15200
rect 23320 14200 23700 14800
rect 24200 14200 24580 14800
rect 23320 13810 24580 14200
<< pdiode >>
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
<< ndiode >>
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
<< pdiodec >>
rect 19610 14310 19890 14690
rect 23810 14310 24090 14690
<< ndiodec >>
rect 19610 27010 19890 27390
rect 23810 27010 24090 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 19490 29790 24210 29990
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 18890 15400 24810 15410
rect 18890 13600 18900 15400
rect 19000 15290 24700 15300
rect 19000 13710 19010 15290
rect 19490 15200 20010 15290
rect 23690 15200 24210 15290
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 19490 13710 20010 13810
rect 23690 13710 24210 13810
rect 24690 13710 24700 15290
rect 19000 13700 24700 13710
rect 24800 13600 24810 15400
rect 18890 13590 24810 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 19490 29990
rect 24210 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 15410 19490 29790
rect 19610 27010 19890 27390
rect 20010 15410 23690 27790
rect 23810 27010 24090 27390
rect 24210 15410 25280 29790
rect 18220 13590 18880 15410
rect 18880 13590 18890 15410
rect 19010 15200 19490 15290
rect 20010 15200 23690 15290
rect 24210 15200 24690 15290
rect 19010 13810 19120 15200
rect 19120 13810 19490 15200
rect 19610 14310 19890 14690
rect 20010 13810 20380 15200
rect 20380 13810 23320 15200
rect 23320 13810 23690 15200
rect 23810 14310 24090 14690
rect 24210 13810 24580 15200
rect 24580 13810 24690 15200
rect 19010 13710 19490 13810
rect 20010 13710 23690 13810
rect 24210 13710 24690 13810
rect 24810 13590 24820 15410
rect 24820 13590 25280 15410
rect 18220 11610 19490 13590
rect 24210 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 19500 30000
rect 18000 11610 18010 29990
rect 19490 15410 19500 29990
rect 18890 15400 19500 15410
rect 19600 27900 24100 30000
rect 19600 27390 19900 27900
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 18890 13600 18900 15400
rect 19000 15290 19500 15300
rect 19000 13710 19010 15290
rect 19490 13710 19500 15290
rect 19000 13700 19500 13710
rect 19600 14690 19900 27010
rect 20000 27790 23700 27800
rect 20000 15410 20010 27790
rect 23690 15410 23700 27790
rect 20000 15400 23700 15410
rect 23800 27390 24100 27900
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 13600 19900 14310
rect 20000 15290 23700 15300
rect 20000 13710 20010 15290
rect 23690 13710 23700 15290
rect 20000 13700 23700 13710
rect 23800 14690 24100 27010
rect 24200 29990 25500 30000
rect 24200 15410 24210 29990
rect 24200 15400 24810 15410
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 13600 24100 14310
rect 24200 15290 24700 15300
rect 24200 13710 24210 15290
rect 24690 13710 24700 15290
rect 24200 13700 24700 13710
rect 24800 13600 24810 15400
rect 18890 13590 19500 13600
rect 19490 11610 19500 13590
rect 18000 11600 19500 11610
rect 19600 11500 24100 13600
rect 24200 13590 24810 13600
rect 24200 11610 24210 13590
rect 25490 11610 25500 29990
rect 24200 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 19490 29990
rect 19610 27010 19890 27390
rect 19010 13710 19490 15290
rect 20010 20910 23690 27790
rect 23810 27010 24090 27390
rect 19610 14310 19890 14690
rect 20010 13710 23690 15290
rect 24210 20910 25490 29990
rect 23810 14310 24090 14690
rect 24210 13710 24690 15290
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19490 27500 20010 27510
rect 19490 26900 19500 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20010 27500
rect 19490 26890 20010 26900
rect 23690 27500 24210 27510
rect 23690 26900 23700 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24210 27500
rect 23690 26890 24210 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19490 14800 20010 14810
rect 19490 14200 19500 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20010 14800
rect 19490 14190 20010 14200
rect 23690 14800 24210 14810
rect 23690 14200 23700 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24210 14800
rect 23690 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 19490 29990
rect 19490 27790 24210 29990
rect 19490 27510 20010 27790
rect 19610 27010 19890 27390
rect 19490 20910 20010 26890
rect 20010 20910 23690 27790
rect 23690 27510 24210 27790
rect 23810 27010 24090 27390
rect 23690 20910 24210 26890
rect 24210 20910 25490 29990
rect 18010 15290 25490 20690
rect 18010 13710 19010 15290
rect 19010 13710 19490 15290
rect 19490 14810 20010 15290
rect 19610 14310 19890 14690
rect 19490 13710 20010 14190
rect 20010 13710 23690 15290
rect 23690 14810 24210 15290
rect 23810 14310 24090 14690
rect 23690 13710 24210 14190
rect 24210 13710 24690 15290
rect 24690 13710 25490 15290
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19500 27500 20010 27510
rect 19500 26900 19510 27500
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 20000 26900 20010 27500
rect 19500 26890 20010 26900
rect 23700 27500 24210 27510
rect 23700 26900 23710 27500
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 24200 26900 24210 27500
rect 23700 26890 24210 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19500 14800 20010 14810
rect 19500 14200 19510 14800
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 20000 14200 20010 14800
rect 19500 14190 20010 14200
rect 23700 14800 24210 14810
rect 23700 14200 23710 14800
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
rect 24200 14200 24210 14800
rect 23700 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27510 25490 29990
rect 18010 26890 19490 27510
rect 19490 26890 19500 27510
rect 19610 27010 19890 27390
rect 20010 26890 23690 27510
rect 23690 26890 23700 27510
rect 23810 27010 24090 27390
rect 24210 26890 25490 27510
rect 18010 20910 25490 26890
rect 18010 14810 25490 20690
rect 18010 14190 19490 14810
rect 19490 14190 19500 14810
rect 19610 14310 19890 14690
rect 20010 14190 23690 14810
rect 23690 14190 23700 14810
rect 23810 14310 24090 14690
rect 24210 14190 25490 14810
rect 18010 11610 25490 14190
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 19500 27500 20010 27510
rect 19500 26900 19510 27500
rect 20000 26900 20010 27500
rect 19500 26890 20010 26900
rect 23700 27500 24210 27510
rect 23700 26900 23710 27500
rect 24200 26900 24210 27500
rect 23700 26890 24210 26900
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 19500 14800 20010 14810
rect 19500 14200 19510 14800
rect 20000 14200 20010 14800
rect 19500 14190 20010 14200
rect 23700 14800 24210 14810
rect 23700 14200 23710 14800
rect 24200 14200 24210 14800
rect 23700 14190 24210 14200
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 19600 27390 19900 27400
rect 19600 27010 19610 27390
rect 19610 27010 19890 27390
rect 19890 27010 19900 27390
rect 19600 27000 19900 27010
rect 23800 27390 24100 27400
rect 23800 27010 23810 27390
rect 23810 27010 24090 27390
rect 24090 27010 24100 27390
rect 23800 27000 24100 27010
rect 19600 14690 19900 14700
rect 19600 14310 19610 14690
rect 19610 14310 19890 14690
rect 19890 14310 19900 14690
rect 19600 14300 19900 14310
rect 23800 14690 24100 14700
rect 23800 14310 23810 14690
rect 23810 14310 24090 14690
rect 24090 14310 24100 14690
rect 23800 14300 24100 14310
<< metal5 >>
rect 19200 27400 24500 27800
rect 19200 27000 19600 27400
rect 19900 27000 23800 27400
rect 24100 27000 24500 27400
rect 19200 14700 24500 27000
rect 19200 14300 19600 14700
rect 19900 14300 23800 14700
rect 24100 14300 24500 14700
rect 19200 13900 24500 14300
<< labels >>
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
<< end >>
