magic
tech sky130A
timestamp 1679064228
<< nwell >>
rect 21100 13700 22600 15400
<< pwell >>
rect 18000 15400 25500 30000
rect 18000 13700 21100 15400
rect 22600 13700 25500 15400
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 21450 27650 22250 27660
rect 21450 26740 22250 26750
rect 20980 15500 22720 15510
rect 20980 13600 21000 15500
rect 22700 13600 22720 15500
rect 20980 13590 22720 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 21200 13810 21220 15300
rect 21530 14850 22170 14860
rect 21530 14150 21550 14850
rect 22150 14150 22170 14850
rect 21530 14140 22170 14150
rect 22480 13810 22500 15300
rect 21200 13800 22500 13810
<< psubdiffcont >>
rect 18220 27660 25280 29790
rect 18220 26740 21450 27660
rect 22250 26740 25280 27660
rect 18220 15510 25280 26740
rect 18220 13590 20980 15510
rect 22720 13590 25280 15510
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 21220 14860 22480 15300
rect 21220 14140 21530 14860
rect 22170 14140 22480 14860
rect 21220 13810 22480 14140
<< pdiode >>
rect 21550 14690 22150 14850
rect 21550 14310 21710 14690
rect 21990 14310 22150 14690
rect 21550 14150 22150 14310
<< ndiode >>
rect 21550 27390 22150 27550
rect 21550 27010 21710 27390
rect 21990 27010 22150 27390
rect 21550 26850 22150 27010
<< pdiodec >>
rect 21710 14310 21990 14690
<< ndiodec >>
rect 21710 27010 21990 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 21440 29790 22260 29990
rect 21450 27500 22250 27660
rect 21450 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22250 27500
rect 21450 26740 22250 26900
rect 20990 15500 22710 15510
rect 20990 13600 21000 15500
rect 21100 15390 22600 15400
rect 21100 13710 21110 15390
rect 21440 15300 22260 15390
rect 21530 14800 22170 14860
rect 21530 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22170 14800
rect 21530 14140 22170 14200
rect 21440 13710 22260 13810
rect 22590 13710 22600 15390
rect 21100 13700 22600 13710
rect 22700 13600 22710 15500
rect 20990 13590 22710 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 21440 29990
rect 22260 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 15510 21440 29790
rect 21710 27010 21990 27390
rect 22260 15510 25280 29790
rect 18220 13590 20980 15510
rect 20980 13590 20990 15510
rect 21110 15300 21440 15390
rect 22260 15300 22590 15390
rect 21110 13810 21220 15300
rect 21220 13810 21440 15300
rect 21710 14310 21990 14690
rect 22260 13810 22480 15300
rect 22480 13810 22590 15300
rect 21110 13710 21440 13810
rect 22260 13710 22590 13810
rect 22710 13590 22720 15510
rect 22720 13590 25280 15510
rect 18220 11610 21440 13590
rect 22260 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 21450 30000
rect 18000 11610 18010 29990
rect 21440 15510 21450 29990
rect 20990 15500 21450 15510
rect 21550 27540 22150 30000
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 20990 13600 21000 15500
rect 21100 15390 21450 15400
rect 21100 13710 21110 15390
rect 21440 13710 21450 15390
rect 21100 13700 21450 13710
rect 21550 14840 22150 26860
rect 22250 29990 25500 30000
rect 22250 15510 22260 29990
rect 22250 15500 22710 15510
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 20990 13590 21450 13600
rect 21440 11610 21450 13590
rect 18000 11600 21450 11610
rect 21550 11500 22150 14160
rect 22250 15390 22600 15400
rect 22250 13710 22260 15390
rect 22590 13710 22600 15390
rect 22250 13700 22600 13710
rect 22700 13600 22710 15500
rect 22250 13590 22710 13600
rect 22250 11610 22260 13590
rect 25490 11610 25500 29990
rect 22250 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 21440 29990
rect 21560 27390 22140 27540
rect 21560 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22140 27390
rect 21560 26860 22140 27010
rect 21110 13710 21440 15390
rect 22260 20910 25490 29990
rect 21560 14690 22140 14840
rect 21560 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22140 14690
rect 21560 14160 22140 14310
rect 22260 13710 22590 15390
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21440 27650 22260 27660
rect 21440 26750 21450 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21440 26740 22260 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21440 14950 22260 14960
rect 21440 14050 21450 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21440 14040 22260 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 21440 29990
rect 21440 27660 22260 29990
rect 21560 26860 22140 27540
rect 21440 20910 22260 26740
rect 22260 20910 25490 29990
rect 18010 15390 25490 20690
rect 18010 13710 21110 15390
rect 21110 13710 21440 15390
rect 21440 14960 22260 15390
rect 21560 14160 22140 14840
rect 21440 13710 22260 14040
rect 22260 13710 22590 15390
rect 22590 13710 25490 15390
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27660 25490 29990
rect 18010 26740 21440 27660
rect 21440 26740 21450 27660
rect 21560 26860 22140 27540
rect 22260 26740 25490 27660
rect 18010 20910 25490 26740
rect 18010 14960 25490 20690
rect 18010 14040 21440 14960
rect 21440 14040 21450 14960
rect 21560 14160 22140 14840
rect 22260 14040 25490 14960
rect 18010 11610 25490 14040
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21450 27650 22260 27660
rect 21450 26750 21460 27650
rect 22250 26750 22260 27650
rect 21450 26740 22260 26750
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21450 14950 22260 14960
rect 21450 14050 21460 14950
rect 22250 14050 22260 14950
rect 21450 14040 22260 14050
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 21550 27540 22150 27550
rect 21550 26860 21560 27540
rect 21560 26860 22140 27540
rect 22140 26860 22150 27540
rect 21550 26850 22150 26860
rect 21550 14840 22150 14850
rect 21550 14160 21560 14840
rect 21560 14160 22140 14840
rect 22140 14160 22150 14840
rect 21550 14150 22150 14160
<< metal5 >>
rect 19200 27550 24500 27800
rect 19200 26850 21550 27550
rect 22150 26850 24500 27550
rect 19200 14850 24500 26850
rect 19200 14150 21550 14850
rect 22150 14150 24500 14850
rect 19200 13900 24500 14150
<< labels >>
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
<< end >>
