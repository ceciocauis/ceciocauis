magic
tech sky130A
timestamp 1679056719
<< nwell >>
rect 21100 13700 22600 15300
<< pwell >>
rect 18000 15300 25500 30000
rect 18000 13700 21100 15300
rect 22600 13700 25500 15300
rect 18000 10000 25500 13700
<< psubdiff >>
rect 18200 29790 25300 29800
rect 18200 10210 18220 29790
rect 21280 27800 22420 27810
rect 21280 26600 21300 27800
rect 22400 26600 22420 27800
rect 21280 26590 22420 26600
rect 20980 15400 22720 15410
rect 20980 13600 21000 15400
rect 22700 13600 22720 15400
rect 20980 13590 22720 13600
rect 25280 10210 25300 29790
rect 18200 10200 25300 10210
<< nsubdiff >>
rect 21200 13810 21220 15200
rect 21380 15000 22320 15010
rect 21380 14000 21400 15000
rect 22300 14000 22320 15000
rect 21380 13990 22320 14000
rect 22480 13810 22500 15200
rect 21200 13800 22500 13810
<< psubdiffcont >>
rect 18220 27810 25280 29790
rect 18220 26590 21280 27810
rect 22420 26590 25280 27810
rect 18220 15410 25280 26590
rect 18220 13590 20980 15410
rect 22720 13590 25280 15410
rect 18220 10210 25280 13590
<< nsubdiffcont >>
rect 21220 15010 22480 15200
rect 21220 13990 21380 15010
rect 22320 13990 22480 15010
rect 21220 13810 22480 13990
<< pdiode >>
rect 21400 14690 22300 15000
rect 21400 14310 21710 14690
rect 21990 14310 22300 14690
rect 21400 14000 22300 14310
<< ndiode >>
rect 21400 27390 22300 27700
rect 21400 27010 21710 27390
rect 21990 27010 22300 27390
rect 21400 26700 22300 27010
<< pdiodec >>
rect 21710 14310 21990 14690
<< ndiodec >>
rect 21710 27010 21990 27390
<< locali >>
rect 18000 29990 25500 30000
rect 18000 11610 18010 29990
rect 21290 29790 22410 29990
rect 21290 27500 22410 27810
rect 21290 26900 21600 27500
rect 21700 27390 22000 27400
rect 21700 27010 21710 27390
rect 21990 27010 22000 27390
rect 21700 27000 22000 27010
rect 22100 26900 22410 27500
rect 21290 26590 22410 26900
rect 20990 15400 22710 15410
rect 20990 13600 21000 15400
rect 21100 15290 22600 15300
rect 21100 13710 21110 15290
rect 21290 15200 22410 15290
rect 21380 14800 22320 15010
rect 21380 14200 21600 14800
rect 21700 14690 22000 14700
rect 21700 14310 21710 14690
rect 21990 14310 22000 14690
rect 21700 14300 22000 14310
rect 22100 14200 22320 14800
rect 21380 13990 22320 14200
rect 21290 13710 22410 13810
rect 22590 13710 22600 15290
rect 21100 13700 22600 13710
rect 22700 13600 22710 15400
rect 20990 13590 22710 13600
rect 25490 11610 25500 29990
rect 18000 10210 18220 11610
rect 25280 10210 25500 11610
rect 18000 10000 25500 10210
<< viali >>
rect 18010 29790 21290 29990
rect 22410 29790 25490 29990
rect 18010 11610 18220 29790
rect 18220 27810 21290 29790
rect 22410 27810 25280 29790
rect 18220 26590 21280 27810
rect 21280 26590 21290 27810
rect 21710 27010 21990 27390
rect 22410 26590 22420 27810
rect 22420 26590 25280 27810
rect 18220 15410 21290 26590
rect 22410 15410 25280 26590
rect 18220 13590 20980 15410
rect 20980 13590 20990 15410
rect 21110 15200 21290 15290
rect 22410 15200 22590 15290
rect 21110 13810 21220 15200
rect 21220 13810 21290 15200
rect 21710 14310 21990 14690
rect 22410 13810 22480 15200
rect 22480 13810 22590 15200
rect 21110 13710 21290 13810
rect 22410 13710 22590 13810
rect 22710 13590 22720 15410
rect 22720 13590 25280 15410
rect 18220 11610 21290 13590
rect 22410 11610 25280 13590
rect 25280 11610 25490 29790
<< metal1 >>
rect 18000 29990 21300 30000
rect 18000 11610 18010 29990
rect 21290 15410 21300 29990
rect 20990 15400 21300 15410
rect 21400 27690 22300 30000
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 20990 13600 21000 15400
rect 21100 15290 21300 15300
rect 21100 13710 21110 15290
rect 21290 13710 21300 15290
rect 21100 13700 21300 13710
rect 21400 14990 22300 26710
rect 22400 29990 25500 30000
rect 22400 15410 22410 29990
rect 22400 15400 22710 15410
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 20990 13590 21300 13600
rect 21290 11610 21300 13590
rect 18000 11600 21300 11610
rect 21400 11500 22300 14010
rect 22400 15290 22600 15300
rect 22400 13710 22410 15290
rect 22590 13710 22600 15290
rect 22400 13700 22600 13710
rect 22700 13600 22710 15400
rect 22400 13590 22710 13600
rect 22400 11610 22410 13590
rect 25490 11610 25500 29990
rect 22400 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via1 >>
rect 18010 20910 21290 29990
rect 21410 27390 22290 27690
rect 21410 27010 21710 27390
rect 21710 27010 21990 27390
rect 21990 27010 22290 27390
rect 21410 26710 22290 27010
rect 21110 13710 21290 15290
rect 22410 20910 25490 29990
rect 21410 14690 22290 14990
rect 21410 14310 21710 14690
rect 21710 14310 21990 14690
rect 21990 14310 22290 14690
rect 21410 14010 22290 14310
rect 22410 13710 22590 15290
rect 18010 10010 25490 11490
<< metal2 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21290 27800 22410 27810
rect 21290 26600 21300 27800
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 22400 26600 22410 27800
rect 21290 26590 22410 26600
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via2 >>
rect 18010 20910 21290 29990
rect 21290 27810 22410 29990
rect 21410 26710 22290 27690
rect 21290 20910 22410 26590
rect 22410 20910 25490 29990
rect 18010 15290 25490 20690
rect 18010 13710 21110 15290
rect 21110 13710 21290 15290
rect 21290 15110 22410 15290
rect 21410 14010 22290 14990
rect 21290 13710 22410 13890
rect 22410 13710 22590 15290
rect 22590 13710 25490 15290
rect 18010 11610 25490 13710
rect 18010 10010 25490 11490
<< metal3 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21290 27800 22410 27810
rect 21290 26610 21300 27800
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 22400 26610 22410 27800
rect 21290 26600 22410 26610
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via3 >>
rect 18010 27810 25490 29990
rect 18010 26590 21290 27810
rect 21410 26710 22290 27690
rect 21290 26590 22410 26600
rect 22410 26590 25490 27810
rect 18010 20910 25490 26590
rect 18010 15110 25490 20690
rect 18010 13890 21290 15110
rect 21410 14010 22290 14990
rect 22410 13890 25490 15110
rect 18010 11610 25490 13890
rect 18010 10010 25490 11490
<< metal4 >>
rect 18000 29990 25500 30000
rect 18000 20910 18010 29990
rect 21290 27800 22410 27810
rect 21290 26610 21300 27800
rect 22400 26610 22410 27800
rect 21290 26600 22410 26610
rect 25490 20910 25500 29990
rect 18000 20900 25500 20910
rect 18000 20690 25500 20700
rect 18000 11610 18010 20690
rect 21290 15100 22410 15110
rect 21290 13900 21300 15100
rect 22400 13900 22410 15100
rect 21290 13890 22410 13900
rect 25490 11610 25500 20690
rect 18000 11600 25500 11610
rect 18000 11490 25500 11500
rect 18000 10010 18010 11490
rect 25490 10010 25500 11490
rect 18000 10000 25500 10010
<< via4 >>
rect 21400 27690 22300 27700
rect 21400 26710 21410 27690
rect 21410 26710 22290 27690
rect 22290 26710 22300 27690
rect 21400 26700 22300 26710
rect 21400 14990 22300 15000
rect 21400 14010 21410 14990
rect 21410 14010 22290 14990
rect 22290 14010 22300 14990
rect 21400 14000 22300 14010
<< metal5 >>
rect 19200 27700 24500 27800
rect 19200 26700 21400 27700
rect 22300 26700 24500 27700
rect 19200 15000 24500 26700
rect 19200 14000 21400 15000
rect 22300 14000 24500 15000
rect 19200 13900 24500 14000
<< labels >>
flabel metal5 19200 13900 24500 27800 0 FreeMono 5600 0 0 0 in
flabel metal4 18000 15100 25500 17300 0 FreeMono 5600 0 0 0 vdd
flabel metal4 18000 24400 25500 26600 0 FreeMono 5600 0 0 0 vss
<< end >>
