magic
tech sky130A
timestamp 1679141029
<< pwell >>
rect 28300 16100 30300 36100
<< locali >>
rect 28300 16100 30300 36100
<< metal1 >>
rect 28300 17700 30300 36100
<< metal2 >>
rect 28300 27000 30300 36100
<< metal3 >>
rect 28300 27000 30300 36100
<< metal4 >>
rect 28300 27000 30300 36100
<< end >>
