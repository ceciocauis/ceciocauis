magic
tech sky130A
magscale 1 2
timestamp 1675091164
<< metal5 >>
rect -1000000 200 1000000 257
rect -1000000 -257 1000000 -200
<< rm5 >>
rect -1000000 -200 1000000 200
<< properties >>
string gencell sky130_fd_pr__res_generic_m5
string library sky130
string parameters w 10000.0 l 2.0 m 1 nx 1 wmin 1.60 lmin 1.60 rho 0.029 val 5.8u dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
