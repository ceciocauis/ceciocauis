magic
tech sky130A
timestamp 1679140823
<< pwell >>
rect 28300 16100 28800 36100
<< locali >>
rect 28300 16100 28800 36100
<< metal1 >>
rect 28300 17700 28800 36100
<< metal2 >>
rect 28300 27000 28800 36100
<< metal3 >>
rect 28300 27000 28800 36100
<< metal4 >>
rect 28300 27000 28800 36100
<< end >>
